��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n�2uO#)�Y>�P[!W�n)6����o�hY[�ܾʰ��)�q�3����ϺeK�^)p��Hz�{%,rU���_��^�^ۜ���l��1An"3�"�����o��LV�laD=tp8F�=�}A1��=1�<��xr7�n�?��;�MHc ��c��Ɨc�ɍ|�w1�ag�j�J�gDBʚ��n�N���a�� Zs��Gb��'�[����_��.#�2��*���|�PNž�0t��'�֩�X~!���i0��A��-�xI'O:1�T���v��W�r�� u���ڍ3�����G����Lֿ�^PQě��zg�nJ����*��EV�I�����u�杇�e,[��l��9Љ�`u6���4�
R�ox�uT\)F�^a�¦/��`ɁK�<��]Ñ�tt�GGe��[�]GO���Ŵ_Kb��f�Ok�i�(���\�,��br;ғD����1�Q������$7�N�����S?L��:�sJ}��%oy��������3�ڴ`��?�le�9��<m�P�y�!�!��sN�E��k�+h�602y�n�AtW�����V��N�"{�042'3����L��l�d���E�3�����Li�&3�����o�����Kk��:h�A�,:qoB�qU�g/�_a1hl���vo�$v����3��4�?-N[����w ���nG2ڻfod�<m�)�������h�x���n.��q��R��^�w5��76�� �8�m<�.U�@�:���i���jH��Ex�Ю���N����.�5p�V�l^�������Ft=֧@{�k;Ee�y�դ��K��Y%��b�ĸA;�QC:��������F��c�A��д�~I��O�,kL�S���q�eH�R����܅�g�2ۺW�M���?�!���;��b��\v|�d����^^�Ȱ�[��r;�e�WN��b���t�w���KĬ��O�y���-�gYդ����m�3�Fbպ����u�@�TE����Ȳ��#���I�>Dں�GgQ�`(��	� `������H�p���X��X��i9p�s��jCLa�'rg�_���ZǪ@��fͨ-�����Ia�a�i[�73����$��.�5��Y�׼2��KÒ�y����$��\�M�/�s��s��4�37��Q�%z�O;h�T_cD~�?���&���YfC��U�PJ.�?	�A�#���dm/�3G��Z7�o/!'ϐ1㘝g��,�P�t��K���w7րX�ȼ�~�����*���bQucv�����H��������:4�O8f9�<̠f]E}�.�̏4���B���;��H��ɫ�p��˭]�����'�eKR����E�"DQ8*�«���¼���+�ߖjv������V��hI/Q��ի��O�=�w��*}���q��Cq��IKL3��p����K!���d���iX#PP�Ź��4������������9�;v�����
'��?�7z�VD-�V'Z&��$���ג��V��5�x�Abl��/�ˣB���uT��j9�*:B`:�#'����-'��V�)���s�J������x.�����Ob�Kns�zX��R��;G3��+?i4(([�w2,�ߘ݅s}]�`(�y�\k��빷�o�-�ar-U���/{�2A��=[�<�(�z�!�lJ��f�v��\CO�١�6!Oj[rP�x
$����f��~k��H�Pp6���Yn@�6�HE�r��k��6d(����~T��
 J�/༚�0nYI�Z��TVR���M4�����XR�)�)�"�싿%Vש��퀷&�CrJ���d
#��0�������km���V���2v3>�$б|����9^�~:�]^k���̀J�0ܺ�l]�8Wp:�4wl�L���.h�e��F����g]Ļ�j��	%���J�x�����6S�t�E�t_�/P�F�Ӎ!4���pA�-�|⋚� �c/f��V�4�����a�W����[,R�J���NY���(�r�wɨ��a ���W��sA;�HB��b��`���һo�E��׊PleE���e�H�];k�
�T������*���Uwd�=�����:�������.j:U7z$�U{���$�w���2��GgF����<�=�#��3ׄ��-OY�|�) ��.4f�]�'\K���#���A�.y(��B��k&�l̎���+=�i�W�7�s�����ib�#�rs�\Q�ٮ�*����� �|b-lbLC�á�3g��{N˸��
80�b��SO����,�g�z̎Ltj�Ut��\_4A���u4ٌ�Q�H�_A_L��T�Q[�(=���m�+�Ier��?TjH����~Vf�S˽N�[�	�N������%�d��]"���h?{	����ZM�JQ��3��Ut�#� ��Y�|��pf�5���Wۈ|pNؙ:�;ԩ��G�4���{8�(�O\s�2#r��㧺���gk�bĵ7�@^��ih�wV�+����U�̚7��:sWr�$#L�w�nPY�$T{����w�rB��$��>�Ur��H7����"���[�C2��,�yd֯e9մ��j2�W)�,e�gfyw�ё�Mt��x�K�.��`npg�}�G=Ш.���k�y��'��R�g����'S՜�R.*tY`s�֕�Na��_$��B%�Dz�5�(�8�"��A�5�t�z�{�|�p}-;ʠ�8G#���LZ~Y�ЬQ���J��Z�\���VƆ ~}�T��!����a|�=���y�clv�����,�@Z��O��Ļ�"B`�$���
�]h,xW~.v�.=C���\��\��׀n������-:ڧ!6��s�]��X�ë<�q1���4��E�g�N'�7��jf��|����] ŷ�geq���*>eU�l��i�=Ig�`���K��+��}	���\f�����bBR���t��pH��;ً�lt�p�� }�ݵ\$�|X7��^jo���Q��%�I��i���cĳ�$ԅ��=-.�vU1�K���X|� �y\L 2-'�w;���So��hvkJ�Y�QZ��|tmE���g5����DYy<:B��S��v�5#�Z�;��iz�ԏF�Q�=����@�E��H�se��6���lh<�4��w�Yg����i���^Iye�j	P"��eJ�nd��3��둞L1�v)̑�_?'��L��;�%�R��
Y(۷D��.>-R����T�����"ۅ�r�Dc<Gv�x�{A9��E���Ro<V�y���X�G�N�4t��s�
��zFn,NQ�If�`�_��ӏ*�6�TIR�U�8$�Iɠ��;p���,�C���>��=N;c��M��A)!e���(�bos ��pz�S�rX�yRfA��6��`�8�(����K��=ց�'�~LC�M&��pN���D8P`~J
A�&�QDIovw��G�c�Ӊ-9�O���&��\�v�빂������9vy�&�~�5i�>�*ߖ��zj~����c��ep���k,���ܠ��� n/<@��k�%��~9�l\��B���d�5�
`O�D$��_R��5O.���R�aa����@��s���ȶH�JΊZ~&��a���/p	��xR�o�Nk��SO�(��j��s`�\:�g�����f��2��^y�������aEhؓ,V5N�zW���X��*��>�\,.�����Q��3Q�ͫ�h��T��`̏r%/���Q7�7�xb��"�Vn��]o�_ ��JXڇ�D�����5��P�zi!�4�zR8�+Æ����`G)�f����S�~��E�vc358ӑ�|C̊���2����6_V������W^i�ܾM�&���r�͑&i%d�@(����.Y;:p�8��vuS�fft�˾Qt�{|'��uq7R��"��6X�!sB�6�����U�IJ!��]���~o���W|��."�DQ�q�ߣ��Ã�WR[5Э���Bv��F	)L�uH��]R�7�<�u�׬�Hj�l_��^�DW��)Ϯ2T�j$ӡ�W�$�R�s��g�����u�W/��	�P�|0�.˽`��3�����$��q�4��&�jMU�{
�n،��H�Ho�5���} 7� =���`����g�3�����[b����v�S� �FmD�9��4�T��=I�dmHz���0���.V�͑�Ü>�>��S	�/����`�9�z�)yM���%j�â rp.!
�J��|l�c�)+���<떊�Ɓc��`ݓ� �������*Mz8-���� �ul S��P�ӓ�ۊ"�ƀ0�!�"�+N�������Haw�zd�DXά�C𒙌���R���ʢCC��\W�� Yӗ�F#�5�ȵ��/��@T?���,sٓ|����k��" ��G��G��F���N��C�?h]3�B�v��4N2���E��}q�|�R��PG���~%)m���#F�kT�*�#/u����?�H9��=��� �����9���ꦐǵ}����ϕ�54@m��2{F��$B�E/Σ��tR���z=�8e���)w?�	V�.�C���aI9Ja�����>�N5����o{W���yw�IlF8qZTʟ��(c
g.�>섮�P�}�paw2YXt5q��T�l�kni#��zq�s�M�>�4�ŚX�,�r��c�=W�Fe�3,5��fx�R�����CXͪ�X��Gp;�G�}���	d�ᝋ�:S��3 �N�ro�F���W�TU$�_}��t��b$P��Mx�6�9��b�� �+��Vt��I�^bw�&-$h��Z���aj�`ƙm�(�����cO�Ǝ�T`ʉͨ��}��.k�BP�Cd�vH���01czǞ�59������8;g�����Q�フj4�����π�{��!�3�B�,�釉%��&)��vY��E+��S$�J4N��"ӱE��7�;��K��>K	*KO�c�����7�	��RT���IN죑#zί�=�"�;�$�U�l3�MI�eʥ)M��T$�!z�o#(�i�w��4siMK�P�S��Y��-���2���Z�y.����U�
>���4����������V�ތp��;1�C�����<ڒ*�����,��m�@��s3ݓCL��� B�&��W�S`1� �
�4�2�oO�V�I,�
���W�5�o�MGH�x������u����	'`0yY�u�]6����4X����]�Z��,�!�C���p����ͪ�	���3�V)�5�5�Y"?t>��4h�Hq%��F��yi����p�Eϸ�*�P�=:�.�.)�o(���
lbn<)�]���	��p!9����䵠��.0�+��t����+	%���W��0d"-�fr�G	��*���ܩj���)_�|%���H��]�%z,��Ug�g�:��#��<v׳���/���|	�߁	�����$1�|ᬺ�K`lߜ���,�:�Z���oSr5]U���j��Z
�W�h2})dk���'�ׅ�,�ȚA ��u�e�K9�h1�I�$��.�`�pI����?�U���;��gk�èz�ui����PW�S��j耠��<���b7/7Ӥ[��d"o����r/>��,k3���'�(���z,蔉� $+�Z��q^�	���Za����A3�s�?��%�|�7l�[�m9��`�TR�r��ߌ�s��t"�]5�/��`c���!&�À4�t��1$A03Β�J�<�G-8��R�F �Fؙ>H�=�ŞE�T���z�{��y�*�_�g�g��i'�!��F��d��k��g� ��A"����=<AE�8�-ef��p���I�4����lU��J����ʗۃ,w���F�m8��i(7��O�g��@���6o9ZT?9�q������i���ԭ�T�8S��2L�#���+W�����c
)�|���w�D��C�[ut÷�"��l�z�n$���q�呶b��9��<��]&��<a���[{N��$�e'���9Tb|��`j�gi䨔̑}�>���E��1��&��v�*�T�D�-흤��@.���9�U��ҭƪās��8[�4c�Y)���	+s�N|M�Y����T��5N�������a����_qyZP��z4ϲ�=��,�f �WkK���ߠ��w�J�n	����" ݛ���e�T�@iD��+O�!bK�-a�8�����߱�����-�?V�x���(��M��眬��+;!�	8}�kB,C��R5fA��Z+���	�J�ks��Z�4�R��n���%���L�nO�*]=@��A�t��X�7����ߊ>*ٜ�3]�����/�%���J� <����F}��\J��A��?���]��'�O�`O��,� ��|d����Us�L�U�y_��ja�zY�
����磧�P�`���	���iɉ�pKr I�,҂~���l���_���u#$��Op��U�Xh��^k��B��筃�t��:�Ky$�q��	�:�k �u
��;T�ي(��Ck;�S3>a�7�md��#;H2�~><��Tk��{�qfU�X G�_��k��K�^z��p�qe	�3�h��7�ҽ�@)����*�Y�&��nŇL%B��`bh~�'�K�#Vȯu�H����!F�5�jG�%M4Ĥ�W�p����j�
̺�sq^�}����B��a��~l�N;�.�@;���jG�6wbO*���h6�`�X9�Ŗ/Ud�]��j���5������F����H]��;�ɜy��XE�%������lt��;A���1ʿv�bolP�W����ݍ�u�>M�B���c��Y�z�؈�����'�K�]ҏR<�bŞ1`u�}�!�=K�V��y	b62۪J����]n�C!i���\�?��a����5�N_Ϊ��Ӭ�g��?]3�ǱsC%��s(��.�PX����� ��}.^��:M7E!NJ��6�f���zN���O��Lc�5mi�6Fn�8�7dUh���+�7�`%6����A#/.h益�TK�LN`�$���_1�S?��U��kK54ၒ�t���`��� r�N�Ѱ����X�A���\;�f@���r�Y��n]+��k�M!�!��`D�x�Y��6�m����ѝ�줼m>��Y�`�4���E$x\^,��\���&�y�x�#	K���z���W��Ћ����<���Ĺ~�$�͵�l�c!H�^'��_�3v�KF\��bm
y�~ߍ��S�Y�	�S�y�Bi����oT��AbU-�Z;�d2zir ��?M̚���*	6�1c�~D0�t���J��'.��[L��I��(���߿.�(�������Ow�%`Y�`*��ւ�t�iy?n��ENMT�rdu �<Tܠ>u��u2	K��'Xu?0���Ǌ���}I�?g����׊��*� �ݸ��_^�z�j^!,0�\�QǭIU���@:� ����t���!Ҭ����x�V��'3��Դ��溡:�"�U������ck���_�-V�	#���"C�@��E$�2vj.�����9	-��N(l�v_��`3��MyON�o����Ja;��Tc���4yW;<�0(q��f���U����;LU�a�"�?k����A�� �x)��43�J����>��i���p�rϧ�i�g��+�	�0��D�� ��o �g�y�?�^Z�ؖ��Z-ƽ�jj�p�tI�/�w�g�o-W����c�ip�y�"c��H-\������Tj�����,b�������	X�B@4�㞆[ɫ�)�ʚ�/F��*������OHY-7�8|��^n�j��܁�����(�?�i|U�1�����U�Ii��]X������RU�k\ߊ�p�_�k�Z}�e��^;-6�7(��_���!��j���3p�_!0��usH�N�c߅�Tn���#LL�Z�e�<�t��F���FӬ�@$�V��Ӈ�SYI���%]�I[�-8�k�"���HJ&����&)5d �Z��= �՘�y#8�,�#�������^�V���3����
��急�c�]f��Ů�iB (���G�Z��xp��P^%|thK]�Uh���.����\؊�D�������C]y����0Xd�$}2k�GB�^ H�|�Ϋ Q�K��g�/���+YOX�jU�J-s5���sETkCi	�C��;�|79=�)n8�Һ�����=�,��!?У��H_�c�@��"�n�Rf!��*�@�FAW�Ѱ8����G�^�Oi+++�k�H��!��%�����$Ĳ�ᡮݢ;[=��D�r36R�����`5���T�w����q��*IWEX�e�V���NT���M�kž&���n=m��+Aw�W"��\n��13�)�(����T k|��}H���2�@��c��Ts�S]:�n}E^E.�i�3���T�#�T���^�u��.����[��wO�t�dy*)\���/�+`���k�ǒ�4j�cO�%3qs4w�	���L�z5��Z6�&��ܲ��-��-Đ�x��M��(�����)�T��pW_tg�����ܑ%�� �]��c��驨%��J��3E:���%aw<L'�|�Ǡƒ�,?��-��+�c�&��͛�n���{�����SD��s��O�>�C��zѰ�T�RԊ�v��G>��lq�=XSU��Sa�`j���9�LRo�6x?�>8���9�&sC���7�!�5W �����E�%&mO�����֌m��>Sm�1�Ǐ��/35���_�5&�,w�3�D+r$;Vpޕ�Y.��#Xa�k��}��=�~Bh%HQ
��A/�P�5�q��-�6���A��uȮ��J�<1;	1��}iT���[��T���H����I�"H��6{\�:A��%��qF�yqY�Ӥ/Ɏ�����D��2[QƦDIy��;}4:A4+0�OI��SL��^+?��ޘp�)$�bΊō:� ��6�b���f��7���ˋ�v��)�w�~�B��)~���$������$x�ac�e�VXE*H�q���Aұ�F0��	����L@E�^�C��qf�סB�R�	M�O�{�n2�lp��Òш�Mb@��[eIp{#�e��^�<󮦓e����+�@��č���?�w�/�.9g���|+�@,�#Z�u��Ɯe�~.}���qʍ9M>��G��6~��@	��H���Ʋ�"f<h#ݦ)d�(��Z�x�~��p*
���S@�e�IPJя�۪ӵ��>m���E��%����Td��>���9��d4�ŉ����_6E7��n0j��"�v�Vi8s2V���:�`�
 �<�gDY�5�8��ˉ����4��Ca����?����?̮�
Tޤ}�!w�K�P��$fCx𖼃6U��L8�~����Y
#���	�7�?�U�W	�=S��N����/�HH�:�vo�} +�5��l����$��|��%�g�;�h��?� �k|����wt�І��\��F�ڔ:�T^v��\s4��F*,>x�V� c��~ɱ9��v5������mMz�yd�_��+uB�F=̶3G�uC���*T��x.|�J�;a���ьь�守<�/)iJM�D#�0Fh�7�%ٽm�+�-^�^�'D.�5�N��iXjb�$>>���\��LqW#x
�2����0V�w�p��G���(r-�J�e���L#.v�Q����T,t"��& �FO�]�K��bۥU~^r{�h�g,D;�O����/���Q{�
C@6�W�U�9e}3`���^D�x߯�+T�[���[���`����	����x��� ��t9g_r�s����:q �r�ѐл�>F61�pƐg�����Xw[�� �&��l2XTqc�k�ͯ4��ĸ�[	ER��(�%�,�\��-H�=�j�I���͘��%�N���@�A�q���F�.6���
�W�ت�t�JPGT��=��� s��:MOx��|��_�V�HG�a5@�������TXS�`q<(�.��S|f�]Z�7�k�1�����Ok�2�t9^g��u��$��#ɩ�|�ـ����w����;#ܽG��[�ѫ��`��a�j��''��ó��_��s�����x��Ů���Twҵ�k��7�y�#�|b��G�����Xn���=��*��}��	�.�'��;2�_n�G���&co�?SԱ�� ���6��@x��G�ֈ����]s�"�мﭧ�v8�wfk�j��#���.\�G�}���pDRN���X��a�A��4`o����5���*ӎ��U�%�U���/h{�yWtG1�%����<��^e�� ;�Q��qՓ�;(tK�
~3��O�Zoń�O��āo�pU���GN����k�mvǝ���PY^f8��Z1�������Ґ/A�CݳGս3�=��j�����j�ƴ���*8��m�K5��`� 2 �*�Z-S�:Mny_�|WcE�����60��^(�*�"5�Ԇ�$fk>sbP��o������3��J@bd�t��
�Kd�"*���O���O�����p�O��SB���3I�F����h�'m<eG���$���YhaB@�3b�w� 6I�;���k/��M��gQ�G'.8�5D���Xkj��M0��LM��N���Y7t><�BI���g	��`x�!�(���B	�*�i���P$jQ���a����o�	zN�ҍ`��kc��E��)�{�������:uC�w]N�+Ԑ��Ձũ�T�
���1l�<_?��Kp�k�޿��}�A����K��q������b��0�����~�=*�88ș���d��p���/q�ŬČ-�aWX����p͆
 ��U�ྦྷ��@M���� T�(���Q��}b�6�`/�R|��J�l���ni�79���1��B%\�BU�禽�qڝ���O�ƨ:��?�%([�*E��"����wE[?��Ѳ X�1�b��~�31U�q�BbJ��b�=L�ԹG�H���Z������u��BG���U[V���ߺ�)V^�۲��УX�!��˫�'���� '��j��߱�����W�b���ejN���)�%UyG���U���*?gQ�֣�\��ڐn#���Z��k�BT�i�&�^��h��PN�Wu;��|L3_�p�Lz�j��!Ot�п���@���Kb�p�����{�	�eFjd�n"�J�?ǭU��ϧ�����n��vVitY�k�����C�f�m"Z�ߚܰ����8�̳���s��@R����XdZx�w�4iL�n^{��)��b�r��v C� �;}㚷�6g��F`_�雭����:ȟ���'���F���4��MV�C��}Č�:Wr�K{�ܷR�����`�<Nf�EE�f��s�%�Ր��_يac<�`g�B��!��v���t�W�{!Sa~�
3���ο�LAfx#+����ޡ���)Z_��I�*<[=�ɲ/�D�I|��3�i�D	4��rDo'��b���D���ՙ�JT�ke �4���-O�+Mㆩ�#(R�O=-��`�L���E��{,ٗ�3ϲ���~<������L��< :D(��B_H.2*�|T!����3�����R�d���c�O>T��-y>?Ȉ&��,ۙ��@?��i��4����Sd,���W�%|�����T�3���צOe�4C�$�`k�	B-%�s���#����$�0,��퐍I��FC�y5{��$���p 	��M�0�Ɓ��P�p���Z?ߢ:z,3�����,�=��Z]��	xԟٖ]��tc����v�jY,Zu�x�\�N`�v�x�y,瘤���Zd�<�80�LW��wm�[�~������� d���Ȉ��iJQ<��za�d�\���X�l|ߌ�b���3z�DIB�8�=� �bV^�P�#�ۆ��k�x3�9卛G��L)b~u�u*a(���� �@Q3���M�i�ҳ�Xc]o~{Z5�����DS�E�Y��^�^p/K(� h@�)	.�&�#�X���)j���$�n�ЧZ��!�g�f�8ŝ�0J�k�:o�}� �˖{�]�	������</�5q�ݶUc�e���ᅰ����y�S���"���e��r�y��d]���;3��ng^;T?'���"$�;���͜f�?p�SnZ�&��Z9�F,�'�k3�؜l�ߜ��:G�l�5���ʱ���"�MO�O����'8�O���0\#�r�5��ɬݠmp�/�6nM��@��2e�3�N�q�^���/��Y+�dZ^{�����Qy��.��T� �sf�#����/�(��&`%��=��/���?$ޒy��Ż[ �<���;*J4�����}D�P�u�)�m���#n���/��C��!R}vy���x%����>;�Iƭ���~S.F�-��y�>z�Nl<e�{���$�����=�K�M��_�y��R,r�ض��If�e���A�Q-䜜�$TH)����NJF�r���w�B.����Ҵ#@(���������~{[�6�Hv$j2�t��ofLXW7�Qh<�qy�`�P���-a��#�Y4v���,���&�2c�s\Y<�Q m�`5���e���-0�h��y@jx���?9m77�+v�
`��֒}R��I:cY�0�	�J�Z��I������Mei#S��\�v�����G�]s]W5�U)�׃��:�N������s6�"oz�*&�vW���J�� ��vq�!\������d�\�@�&��:e���$i����ʃ,O����=��+,912v�������F����aEY�^��8�&᫾�x��e����Hu���a���Y6�P;bHC���aP,˥��I�j����	��ܷM>z����ZI2���ed��	aR��^<���?YIu�#%��j�T�>��ҳ�g�\Z���1k�-�o��B��d�ғ4����4CH2�I�F�d����λ�r��k�q�^
\C8gUu�����z�)���	��`]՘��db}:�O�n!ץ��ջ��]7�ylY��ݻ��Fg�@I}��c�<G�����u�<�,�<UHm ���U���U�Җ7eŘ������ 欂iX���D��"խ�JO(a��~b�%&��	�&�@�1����)�qJ�Q�ڔz�4Q5boƏ��ȍ�^�I7=!=���>���zg�Y�-N��	y�� {V�L�p�
/d#�>-��t���P�h=J�:K$*4�cf��RF����JSn���*��]�(dd�p� #F��$�9p�:�:�F9I2�`H�ջh��[���W������c�
	ɛC7� �+�]�b ��(��s�\�a��2-��0u��)~��or��S��:����P�6z�oL���C)8V��7V�����(��4�h �>���%��8�$�('��[�yʷ0� �%��~��Q	=���������8�XOj���·�n.��>sK��u�lI�
_���"�!23�fO��E Eb9�%�U����z���Il��9Z,/H:����� ����h���Ј��7���b�4|��O��x!	B��Z�>%����F��yu����<=~�Fh��%73�	 ����C����ְ3
�hX�x&x%�Q�l�u�|)'Q~�b1�w ߽m� �Fr�\&	�WD��#	�B^��7�T]w�Z��bIA�Ck�I��<��	_$.�������x�̮)�޳B{`�1���<�z������a�������On�{n&�pѱ���Q~{D����q��z�Y��?���A	J��G��x
��3��������&*|{�ԕG��%���he�˸�-I�Ah���طy��в��A%b��چ��5��;4�%]�b���7a�4j�â�$�,_��M*�1#����ƹӑ�4);����%�B�f,���B�9�>z�J*�(��_�A�[m�����=�)Y�`�*��� qM��6��t�TM��2����fb�	nm{����n�%�٤Ɏ�u�#�����n��vxc�>��#|�M{�[Cѫ����
KM�jZ� �x����M�Q�.k�����;q��_���f�'��'�W�H���A���tC_{�[��iߦM��&�8���K݈k���ja�,��*X�sʇ�*�E��J��?��?�J�Ώ���!��R�{��cC}����#�����Vڎ!0�#�i��U}�e�!���W�5U�<����N�ĪQ=q7�塤EaR�2�̈�ϩB[r��q}�@�S^VʧP�@�
T�+Q	��&�.`-���˟1B/r��8�4pT���Ikkdt$B��#D5�3�R'���V���l;_LNC�aA-�yO�J�E�u�y� �-9�<�k�$K�rW�=3��r�6_�"ޕ���o ��`�3�-���q{1�e��ǝ��4ہd���2���<
�k������Vt^��H"�� ��vp�~���pquy��X�(�|b����M��||_�/\��2Y�U�n�E����).g�����|�w�X�f�s$BzCNIFI�d3m���+�r����XQH�b�;/��W��t�,\OP��F�<�A��et�p.�3@U���~A�b&(����{�s�t���St��V�s�qהL�o�*L��f�T�aq�
d��B�t�oI�����i_u�
�Y��xsB��t�_����O[�����o�c��c~rRg岃���~&�+yH��?�"Au�8�5\i��1�����w�m��ώ�r�������Ag�U�:\�����by�����f~�>���?7FSa�פ�]x7fAh
r�?2-ex>U�7	�Z��q�G�Z�������:�d�Mz��wY�����,7/�+G?�,��݋dV�q49��u{%��e�db���0��V+7I^t�z���v�B����>�2��ǡww���@n�
�!��R�>�!Aט�;2��`=K���� �r�w��g��h���+2�$u0�s��w�h���1���`�{A����W<�?��+�)�e,۬o!%4
���d+W�Z}$�e����<$��d9�ϓ�h&������U";�-��obr���y���L�|�X=kǙ�;����X��@i^s^D��J7�Q�?���aa,Mx:�B��ĩ^כ���C�bu�z�	��k<L�A��-�i)��1���y�]�q��Jf�m`WF4d��Ex
	K����G�8�@l)Kc���|D��&��Je�	R��@�4@ �T7�ӈ0�OkB��Vj�T���_lq�����'Ck�[�N����]�oRm�?��=��3.�Eo�&�Bpe7ǃ,}d�J�Y���,>Uow�߉���0������(%t?�%��)�������o��D]S��T���֔�qG5�!x7���d~��A�E��h�`t�Xu��<�!
���n���_)��90����r�b,Pj21��);e�-r�Y��m`�K�N���T_�kI?E�ԃ�a	��J��� �߾�:�j�_��˻3����#��K³��O�^%���L��	�@��ʽ��Mg�X��|L\W�$کI�($�Db�� �ڞ����>���}8���D
�S�K�g�U�O���̥A�B�tJ)E�:����d�;wV\]���GR�ef%�;�ㆍbH���b݃g�)�dc��b��Y��������3iq���O1*�b�Z�u@�r2~ �9��qϳ�~����M����myd(]�b;�6s�ATg��ra��瀞C}�خ��Q���^���H�}?g��h� `dPЯQh&�w�DY�B����]����t.��fI42��TY!��I�A��O�膻E`Ly��Ԡ��գ�ШC��e�yۜ��_�����j���/����*���gʹD/v�3%e\Ho�{p5�!H!�� ����?Dv�N-?��Vx�p���V���EI��.�]����+_۴;\�e��,��"]U���!J��p=+�J����EE?,@7�@׌��L��賮t
u0��fb���7�	�/�(�A�nٞ��7�]j�C,�Kֹ�	��0�.k��� ѣ��:��\if��:*|Ԧ����f��%7�������7�v9����[^5��ϵ+O�ѷ�h~o��X����2����sB�l3�.���6���O:�U���/w38�v4�^�������a�oN:������s���[%cW>:-p	��p#�ǯ9u��
V;��j尗M�����pH!~�1�R��|��F�gPz1u�	����  �[S�1U/x�����G�2jC9�7o`�!��Q`vo�>���ޯ�i9��'�7���
�1��'Lq�� �i)0����6���W�s�c���tH�:�ϝM�G�F&r;��~Q�ge�I���f����<$W^B^բ���(���Do��)��C��r�(؍���~�J�AQ�fj?���vJ��)& ��rc�$I�㥶픂4����1ue��`�:%���.�U���]�|,9�y�Sp#MP4)��~_u�v��>����� �B:��(5=��  j�u��x휉���6��̥��m���	:��" �t�1kaw�@E�	��K������BQl�)�C�!�>0F�<��46n'Q���oF�J%�O��kW�;U����.��
�!n�)m��V��b���S >\��3���r�s�~�vꦡa�K�4�=fV��y'�p9�E��To �D����-ri�1b��Ձ���eC�|�\�ĠS0dJ��zP1}���e�
µ�A4������xBx�g)G����Lo������������K��N�/�`��R>�h0Ι�ۆ4x�J2G�RI�.����#R��7c�g��evVҬMʈV��2��b�X#��(�8�r�����>8u?�M�6X�G�����8������2\��e0��*D��Z�<Ip�U�iW��:}w�7Ӆ��k��x.E����-����M�ߔ����/M��?�mP{��{=nԒ5x?���uJ�{��������|YO�Yf����]�^oG�#�k�.��5�`M�
�y�ˉ�F"�f�+q�^����$.fW���bT��������s�b	�?�p�Z,H�b��X�NG|�]C3���9=F�t�R�����6���&���X\����cq-T����|��W<��œ�|ۗ4!���	��@K�ň{� o�FG2d<0׏GhAǷw�X����6�o�nԬ�]����?�-
V��!�TOZQ��A�P�qk���36}n�c߸P�s���L�w������f���
����+�5�����C�*�B���� ?�я����ޕ�K���H�ݑz$Ӯc'\o�m�}{����l�4SVjy#	 
�C�1�S���v �y������I3b)�'Oi"�>�8��]�`��*Z����bq,�F8�M�	�c�q�,���_-�q����}9��ͥ!�r_v���vtr��dyA@�z�{ȶ��;�+0�x0���Ӯ^Bq�����w�q��xԀ��N�dԲ��$�?�_9��0ʗ�{��T���5���M"iI.2Ϳ<�о
x���2��c�f+
7x$�7m�-�6��F�	w��Ȟp��-uc���@�%�����2Y8�t��t�~�e���,M[�lN4N*�0�a՟���ef�,����\������T�G+E��.�������w�7�t��z�R���ޛHiYi�����VI�B���1u�����%�q��$[ٞ�7 �}��N�����?�%�m�
�}_��Dr/�q��[��$��5�7�n�\�!x���������j�j��%!yu� �����`�Re�=����Jm��yĄ�!�	��N�ߠɍ��!�B��+�L �Ub�yV �/����E����<�Y�sH��~��ӓm�wj���C��Å��q�)��Qe��/2�{�,'�
K��,��T@Ӹ�D�$ވ�����X9E�;�O�hy*[�5�ȗ B��#Q� "j�~����u���"��ܓ�<mk�$O�)�uv����\�9��>""�Ip�4��f\�����eX���N�A�*���\{1ov?�B ��'fؚ���zl��?��i��7�!�|�rǻsfUF͆��;7����ta震(z��&Q�s�v>a�_�����4�q0����@ї�t#|_QPא�,���r�4�������Ij�l��2��ߥh���U���}���]��TK7���i.�Yw�T�O&Q���[��ν�N����DyB��貎$eL�2��s� �W�o��q�i���\q���`��8k�fe��5a���g`�0̭,��:��~���pB=�ɓ/�w�;����g�$ ��7�Z�[���o�"l�s*��k���`2��W�I��ol�v�{��";����������Bӧ$5�q��ڃ������&���&�T�;!d->}�b�Tc��;�x�#E�lJja�Ni��ܙ��Ŗ�?4�l����z~�|X9�}�^�[Q���3�N{��<�"�#���g��&��u���x`�䑓�qM�����å �ж4(����VK$N��_^��Q�d�^g��"`;���r���t����D�E��}cu�{��F�3��L������s�XBb��������=6�퍡ĕ�X��.������W�ƅ��ՠ/�\Cu�.�1�"a�_�[6��`3��v������"a�/�7�$Õ����l<{|�1ǿI�<�����|��ō��K�v��e��:�Nk?�,9ރYI���F%M�8�L��a_ߏ�`�s
M4�K@d�x���:Cc�i"�
�<O$F���NSq{����^e��{�C֨W�,`u�rp��q�N��A�ۄ���p�b�5ʪ�{I�d����X��,_���~z"��)��b[V��}�4���̂�� ��l[:t�q������T�ϓ@Q^�Y?����<��`j�n�ܸ~Ѩ<>1̻���~*:.��1^�e�# �~��~�C頤ս��pY�)��Z��o��ِ�ԭO��:��x�KW�����@t	
륩��-�M�{�I7�!)�x����'�x�13�Y�_p���$�_���f�Q
J	���B���
 \�|���H| Q�K/"�Ecn҆L6io�sM����|�=n����	h�*n��'�I�$�x5F%�R�
��}�4o�-�nE�C1R�G��1z��j�p֮��[Ǝ�ح���|�$aG���ï�3i�Z���PE�L"԰�'�G�q5�:�OӾ�����n��(!�ƫ�u���/Z7���J@&��vBL��v@����9�!O�i��0���F���F��:�{��
��7��@"4�F���M�r�7�����۫���=��+��+���Z�g�ĩB*��hP��<ku
��Z���Gt�F0Q�|�0Q�EM4;�T�T ���K&`X��^��pw�����Aޙɋ��V�vo!�����Ak�ӱ���aI�/�X�*��(�~������CG<<�ct��!��l��n�@x��������Gz��}��bŏVZ�Q��58��0	��w����s,�Q����S�ĳ��hd�T����ڤ�R�4�r�o���Y�tϞ2F_c�nfh'���cg'>�*L����+��h���l�1X�[� gR����b0�A`ZuA�;���������xY��Y�eãG���9�E�j7Ӊ��2)��l����;�R�x5��ig��?w�Ne%�.�>�~�%:d$NQ�a��p�",(��z���q������L���使�Z����dڬ+��Q�͢{�hK��P��.�$�>���u���q9�^�u/L�Z�"a�-K�G:V-^б���{S%^�;���s�����]�g�,0:�+]řj�p���_�/���+ �*���Lf&�5����ƹ~N�t#���i�o��;��e����K��|<��s���jÃ!ʱ�?��N���N��^�M@>^�L���:�P )���?Uѯ��r�Q���+[�&���$�{��kǁ{ֺ��ۗ��kbzߘj4�%p�U�´����k˺m:?�E!�1��S��/�"_�uE��{>���9?N,$"��Dk����xi�!�Z�6�4������"��z�,v�n��S��"��$��TP��1 }�(��Ea�93C�k�kF��q�*�s�c�{-Q݀�*�_c{�;:h�ު9g?'6���B�����ѕ)ݩV�v*o�0�X;y��\E�[w=QdS�,���(M��S������$����q����i�6��Ҥ@�m�t^dw��g��B���Zx�h��nZ������խ)��,�Z�<�0n�����|��<z�"ӁT�'d�\�{49�Y~�+��&���Z���B��3�-�8H��m��d�ܳҽK�(�F�6���]�����׳����W�b�u=�v8�!8.��&�����a��t�:�M."�܅d8ҵ\�k-����F��m�W���NJ;7%���� �k|���|C�}��ov����y@Џ��L�U�� ��Q���}9$���@MX�h����*���k�AW�ѳ5	�/@���{�����t��o�s��z'�aZ;g����{3Fr�n������֠�cN5,a*�'�&���
.�}*0�x��*��\�$BG�D��1O���XL�C��^t�;��E�~{+�.ߠ�糩��_w��0[K"؉�ꊏ�D�YM���Ɵ�FF޷�$����D�r/,�H��i�s^Eg�-�8�;���nD���-H�j��HYε���(,ώ���C�,��J�j��b.�yUZ���`\kq*��:O���/�DI�1h.\�[NZ����Ӏ���c�nˏ�@����M�KV��ƽ�a_�#jU~�?ڬ6���y��E	M�
���B0��Kh�J���1�kx�@�y��!p�P������Ӈ�S0�De�F/�75ޮ���@����9r� ��:l�xV���f�$q�0M��~�X��gy�:
��	��������Ip�os���9楹~��T����i����{�y�t�;ds�Ip�<�O���ms��|��%�������zz/�>����.9��{���70�ݖj�o륒�G�]tp�j���,���
<A,X�Dh��;�U�����R�o�R~DCc0�_���A�O� �QMt1&�[:��5t6��'��K󘣥]�}a8�76�²F���|­�Y��c��L)�w�~Yl�m�W�f{��ʱC#ffƢ�+��xӛT�'�;.�9�>_�>�1�<�/~�!�ki2���'.㿛4����;pK�T縒�����h��+X�pQ�r��hJq����mܶ�RK~�k߁��F���=�p[Kw�|�|_����[�f"�BǙ���5[�ݥ�����~Z6��9�
��i�_g�X���ѓ��w�+eF��.���s��h~X��7Z�y� ���z5�+����<��dS��I����ݜ����!�D�_��;Uo�xcs���`B�D#�u����a0=k����dj.os�`��6�a�f����P�c��@0h�x>��(�&F��+���������ZeQcm6�ߡR�Z??S���J��VB�B伤��K=��²W��������jʙ3-�\�9����?Q(�A�dv�qgoQV2����!�3�r浛�;�D7�>v���6/�Z�U��uB>bI/�>2�����8��<�b_xg�r���r����J&	�8^Jۛ
���oXmb�Aٽ{�-�f��C�¨��J}�}���681�,5�w��;;o8�D�Gi�5��z�X C��3pg^&�Q>`�ڮ�C���SL�:�䈐Ir��w����1�}��po��������4��=��q�|#閭+�>a;��n�A�"OU�:�Jv4����
mj����@t�}�	>��C)�6�=�s[F���%�h?^��!paᡓA6V���ATU�ga[�P�hDv�������;��c���o�ֻH�)���ۓ�?XK�"�De���<�>b�#���h�a��>��l��3����W����������x���ɻ�lo�J5�C��=��*H�^�F��n�Mud������k.�lF�2�v�<}���^���*��evhܕxc�T���H���Ua3�L+ٳr=��P�ҙ�ԩ.�U�9R��~^����[�ނ������yr��;ݜ�j�����Y�����=�"X��!#O��$:O�"�IpҰ|�z�@�5���}���C�Bq�7���y��$)��!蔛Qc�uc�9]o*����+�vDy���A��s��C⻁�1 /,���u��S����U�r���?�:�T=�E�J^�Y�"�	���`��z�y2��ʴ�$���%m���Φ�t/�]�蜠FE^[��0��z�����&M�wu(Q�9x�#3�W�0�|9d�Uk\�	�ů�W/N1Moj�����<���l<TZ�i�9V��������`��e��E��|�Z���=uR)��^4���\����bL��W/� ͢��\�9���@_������fU�����a<�r�lޖ#ࣹN���xx��]��B�P!���Z�"O���:��&t%�G�����ͤޯ�)|�E�߇e�BK{t�Kx^2wo���`��ck����G�81��JJ��ǝc�����0��f>��#����4`<Do���mTKt:�9�V�#Ru �Nz 3��	�V�5�pP�����ab�G9`G�UUV( �����ţ@����¤K��r��}�ID����w0�(9�:�� 	���9ئ\��451�^D�v(Z�t��x���6�8�F9uY|�K]�N�QDW�e�����鷊a�ys�!ǻ��9b�8�����i�n�f����� �v-I��5��(���l�w�G�)���
�ûl����6�CU�[����L�� N|ֲi��cMɬ�876�t�h��x�d&u'>!JEk�vg�¸�)�����M\�����ʝ5+�pڈ��79�� \E|W��P5�*�X�Py�:�J��5U=����\��5�-�@�c�Jw��,0�֠��&hљ����gĊi���05����؁7?�ە��fY�HҦ�*}����'̕.^��M�� ��]�K1j�� !�_�ç��KX?������t��4b|���YK�c��MW)��1���<�!גB4��U��|�zk"�4x�e�Hy-bo�x0��\�����?\m��so8��Q�3�_��'*���fHr���H����Gt10�M�rk�Ru��,*c�\�B�~,9l}�� �t3��}��gp܀`.�-���儇9b�>Ρ��A�~ґ����\n��?P���u���+�[qܧ<d:�S����-;̼���$��@��S�l���y ���@����.�ڳ����;�70�L3E�V���;/������r�/L1SX�u���{��ɞ�w�tΕo�K�~}��N����Y����r�x�|��i.W��ZL�i:Ϧ^۰��h��K�ǿj���F^��\ƫ��^�����w���ԧ9'X�E�-bp���*t���Re�V;6�z������wk��
�Aʧ�j��f�Yn���Y2͢�R���S��@��7e�R��)�K����y�)�D]�5�:�"M�%��~���':���v?�8FY�	��A	I]��j�,�~��a�m^;�>�JmR>����m�mV�@�KB�E�b%%E��A�u���8�@h
�՗����G��{���M�,!�W?�vᩡ�:K��hh��/So1�lg-ƒ�/�$�`?HY�X<m}?��뚆x2^h�E�¢��d���pX�jN��2W	|�b �Ky[W"�ζ�V����\ULb���CZ��l�[���pr��m7�A⚱'?�ʣ�z`�*bI�}܆z�#�΂�@!��Dv[��*[(a�E��OM����F�5���M@$F܁	�|��MN�KG��s@Z��H^��)W1,%2�6*Z�G�zub�qm���;�=0qd��M�<�N[Y���|W4�}<Eg��#J���gK�q ����Sj�F���_�v����A2;�x�pE6���:4]��~v����U����8=�v�%�Fũ�6��v��a��y!�J#��Fڰ��{E�#c�I����I�6�9R��Z���N��k�mMh���A�
��h��y���a�PfX�����R?��~`������\���$�ۋJ��6�߉?I3vf��!j��1ۛ�@�����%�t͐���/f��dI��V�c��;7B�%�M�"�>��S/�:�]TjTJ?�٤ ��l=������H�-���@/8�����U9Nou�E(ݿ��8�A�?�M+��H����}*���p��X� :���r{�81����<��������b��Ա�7�I%1�tm,��X�[��λE��Y�Ir4��y|�yS���uig�L��-(6�˱�?h�[��T� �k� ?�a!�*��R�.C���Fa��=��c���	H
?=�O�h������s�"�<5b��;�FȐ+պ�lw�7�s�s:�
C���a�&OI��'[�+�\��|ߝ�9����bY��!V�2r�e�T�1�=u:��I�ޗ�~�;�atv4���.��0��z���Z(��Hͺ;j,l�fRF�m}#:*㉐��@��L�>�ϯ<�M��;��d��H|���=	��U�g����if����Ʒ[�9��sZ �FG�c�7��o�(���W�-��(ӱIP4h��:���!�Ŭ��p��ǽxq�߽��N�#�&�Q"��Nh�����11��/%ͷ�+�m�)3a����=L����5<;�fZkm?��I��,��EJ'�
]É"MA0;���d�nab�Śz#���ų�e�$	�����9�X�`^-���gC�U$�7`a�Vr9��=ۀ?b�@���=2:�p��y�8����^!b����s���a�
�2�M﹘�6$ޞ��=Xn!3��D{�+�X�2�����vF�q�{?��R�wnFW�3�J�(�[�=�8�l�bM]ו�zׅ��S�+��R�q`�_H3��[ā�[��PG����h�d��Ī"V�/��p�J_|-��j!M$"�`�6&<���@~y�J�8ǥu��Su��ch��פ�8(�RJ�c��ot��U�Aeiq���*e��\q�q�k�PM������6��g��(f rpr/��D�)G�-ϻ�D�,�ĢqG��)$ޛ��*�¬��Ȓ��wW*�[�j�^)1��4�1"�x�=a���x��� p{
q&s�P.8QҬ�\z	0�W�i5�v�1~ͺ�L� 3��+���yes��u�(�U��
�(G�����@9�s�)���}���9���+�5�L��8��e����Qjy�e_�6(���5��4��j��1y��ݺN>�k:(B�/�%��N��u��*E���������������\�>�]�U�����iCPh��6Q���һ������7^�g�ͽ�{�k���_�\�;YNI���ĳm��l
�ն�Ƃ���*D{e'8����W��p�4)Lr�y�l�Ԯm�-G���,�%�B9��;�Bu�����Z�pt#���:�	�tW�Y�S�w�J������G����+��?}�ՏЍ�_�D�D}|b��7�br��s���3����u���U�Y��-W@�6�����_+���e��7�^�8%���Y�!��et&���#i��0��	�&5/M%���~�SVEb�[���J��b7��U��7�a�탺-_���׻��߶�lV�Y|l���<��v�-['7t��50Vf=ޮ����84<���G��������а{x��.0Ɇ
n�'����H�7Z�ᒯ���t/����4i�T��<���&}дy<��g�֮��!�CfM�頠:h�\h�]�q�P�-Q?��	By��Hk{�1�(��P�^1e���Q�:w+���U"o��#ͫ��5� <*���=�o(�A�-J3�����9�����E/���{Lu�Lׇ�/!e�L����.@�#�⢲����r�􄰘K����$'�Kxۛ}�%�O��Qǳ��ym��1�V�iС�W�B-0����)cI��ؼt=������G�:�6���m��_��Й�tQn:lI��w0�����%�ϣ~�!i���uv4^��a��R�|�:�m�ۦi,�t���D���-�� q*��P�=�h�EKOEZ#���S����+�w!�-~6�L6�"� qI�4����J����1Q}s&pF�X��]l��a��ؿ���MM����U�z^�r(L�XŋC�#{�$J�|�Up����(����ڮ�B�t( �9f�aj�
Щ{Rز�gӁa����#E}K&���']�zg,�8��;��̈́<vm����~m�,
Nd2�s��y$th�r��������{O�x�)O�kL�N�.� �@g�����d����M������0~;ڄrb��PW�4�/��b}��Y8�9�)�v�-�]�G^�̥��\��4��w�f�%���j���s���1�P,<A6:�7�Q���)�B#�R�'N{��y+|����ζ�|�t�����Q�BP�|!�!�q>fz	Dh�#'�3w���e�3sz����� Z$8����t�H�*�Q[�p�&Ι$5��6<�~�t{f|cF�Y��1ᓳ45�����_vمpc���ɔ�����.x�I�g��9���+g,��g���~z���VM���Ǝ~[+U��k"�Ig��r����ZN�-�1�q9�NfE����_}g?XS�Ѩ�;����8�>�|�r��H�� 3�1SL&` ��]�$tS����#��_�+3��w���N�Ey)U���@��A��~+!��[
��x�#��[+�8���	З�U_K 7W���mv��Ȕ� ��1��k�ջ�+�+"-/	�]D�v��%!�{��-�>�b*����p�tw)kpy�����'A�?��vc6��Q���	A��f��M�ǔ<r�t�n'k~�6T��$5�ˊ���ǫ��>)H_����r��H́S�U]�X��� !�r��4��|����i�+�� ��W�Lj�T��R������T��A��+���b�S�pQ�Y�%��aoY�c� w�ovr��}�Wzr���Ԙ���c�U�{0�5g:��[Qݍގ8G��O�Q�k�-�L�R�0�0����?��j�at�\uM�la�Vb���<R��'����6r��|��q�����*9�P=R�a�o~�6Z@m�%#�-'�e�Jd����pT��a�y�W֜��T̹���@=+`0g�
-gLBycQK�[Y9 9�Hw�K��|Sp;zRT��4�@����/��DYro��Lgu�Y35�w"�d�o�T�����u�1�P]��
�-^�O̶_Ut���G��Ƴ/1�)��_�}|&<b�&���*J���
��2�X���&S�ɤ�tC�5f./��m\�r�{dRP\����,�Kf��V%�V��lp����K����;����x�R]*Hvn>a�19:4Q\�7����d�*&k+=�(�x-�)8[_�I����X��űY��D)X���n�"��#��^'n��|剡�7�JM��^���[��ڸ����rd��a�xb�s�VDM�j�E�w7e�R�� ��/4�E��J�l/)kL�f�x��A����T�K>'��v��0�@o��H�o�|=M���Q�u�P���Nm���2J�i,�f��2��^�j��P
Kt������#Q=ݙ��x�@e������eQOQ���c���������l2���^�b��e��Q���,���~�AI��AJ���g����FN ��/F@��Vm.0K'����V�'ɨ6�f��^�Bf]B��4����k+젒���H@&���-���n�i�t�ʯ`*���ئ8޻�}�|�1�G&�܀]�	b�2Q�L"�r�61 ��)�e��A��K�ߋ�\�!g���dm���!x�����Wp��s��F��u���M�)������R��,��s5�/%haij�����P-�v�As|j�Y�P�����|Vd��7�;� �ܞ�da�w$�H\����._1q4�Ir�ُU(W~&�n��c.ˍl���+,)�2�Y�����:�E_\U!��]<E)�@�<�GL��I��X�E�{B16�fa{V�,{�E2��;x�b�9�o���]��3,z�'#��&!w��aR���Ed��:^����K��,��_���b���۔:�h��P`���d� -�hHJ�g�Tw�.� �;5�γK��4�gb���,�\�{�.b�vK���
���ɮع4%$�h��Bu�;%ѐ�q[�%�cw4mk�xZ?^�aC�l�~\#��Jx \��E���9K���6 ��������d��RSӣl�8>����(G���N3�/�t�k�^�:�E����
�6�ª�� %Y�Ǚ�m�NF��`U]��\����B9V?$[JF�7�?�\��u�/t�tb�6N�REe/~d�,������(B+�d$kP,�d���?����B,:69c�wݕ{X^(�K«�B��"��*�\o��Є�v#C����g(JM�4Ha�xeY��a2�l��E�Oи�ߊ>��uq����Mf��ÝL��y�
�H*��h��"� �6�eq,Vkn����^L
w-���-ﳶJ_\KI���	+��%tJP�JokT�.�\y5�_|=����:�s4�Ӊ��ܩG~�ʖQ���I9'�D(z���O� �`$�^Q�2I���k����r��?�Z6|�Յ�M���ͤkx�RWse���X�q�|T;:&�&�L@5�{|"�q��g���^Z��`WY�bv8Yx�<9�����Z�M�9�#��:���cf0M��o�9�V�V��gpp��u�V.���ѓ���L)@��6]#�o���:M��;�{�Y�~��s�I3W�-Vr��U
	�K
C�����k�ތ� xq~�&/�N�$��h^�3�6vx !�/ޟ�fQC$T,����7��x�-��3 �m�x\��Gk�Z��
h��",C"�K��R�od�/h�gP���< �#c_�
��X�B
���uX�x���o;X\�
�s�#���O%����+��K��Ϛ:8qB�}���'uk�$��aM�Wb�gsJ	���x��WK��gì���T{�R�ԝ�K�jt�Z�6��5��;�â�y;��Ič�j����x��0�M� �7���p�ZoÍ��CN5��Û� ��i��T��T�����~U�-�9��}D:�cĳ����էÅG�ti�*��dF<"�	��g(}�\�"�U�Q�"�������9���}��vXe�@�%�7�R�\�<ߒ�C�i.C��@r�(�Bq%��]��'�.u[o��z��fۻ�*�Y!�,';-�D�݄�Vu?���,�,kw�3�ỎC�$yރ���=�q�f��5`2�`^�|��0�f`�aH�`���r��L�p�/�R=�RNafѩ��",�4˪wv��* �S�Y"�
zQum�Ă\acPn�5\	���εεܠ#�/ ��|����V���"\���'�\��iR]}�0��6���R
H"6��⬾�a�(�͒���a}>���;`)���%���|�]�z"@d+
��pPԜ�ȋ�7�4E�i�U�d���c�|@���|�>S������xH�	��&|��
����DAЕ�N�4a>�(�,��C�Oga5������y�*�q�&�S�;s��Ƚ#�Ϗ�n�]CephJH��].a7f~������ ��A)�����<�&�����$�3<Z�|Q*�6�4�3���� 6 <�-w�Ro4�ji)��z��S�X�}U���A��<�c/�S���BA����uu	g�^ܸ6�����[3dP�� ��t�����K-�n3���݌=��J��B�q!�Abq^�N(���z1�T�4���Ct�,�.���>l�5���L�K[�:)��.E �ĉd��*���+J LT��S�����	D6���r�ʧ����o ��qњ��~��/��F��ţ�/ԏ8Ԉ�ܿ���(�U��N�o\8b�s���WWJǶ�(���E�eIC�̉+��ƊU�mH��R��vGC��'K�1�HX���}@��Z~�;\��Z[߻���~6O�Զ�)�x�7�[G僶�Pe�Gs�.gU�`n,��J$Z@�R�n�ΟȀ?�����(# !
��K�vd8x�������$|Nw��5L�ˆ^03-{�
�Z�s4Si�GB���Of8;p�A�f��Yݱ�0V��G��00�9�D��+j��]p��O�v�C���,,��EF�2�$8��6�uu�\�I/?(u���2�;ź4����t(�� �o��)l�WV��͢;n��GF( ������!�j&m��3�9��N�
��ߜ�@��nw|��/�P3p��<~��F}.�u�Ӆ�皞1�W�?Q��pO�qM��մ�!�7#J��� �oG�X��A���B7ej�Ɩ��非d̢�����x_M����E`�TZ<�*jP��Zpz��f�x�D�PW�VI$��S���m�y�A�#E��N��>}i�����El��D�<�wp�&++1^��#$U��� ��ǼQ������U�?ߩ1'��A�o�8�4��;4�C�n�L(�\�������� V��aIn�\Ǳ�]%Jz�Ijc΁܄\.�C ��&P�&√�},�e���t�!�$�.�_�Z�R�\���3(3�oH��©(�Ns��Wy&rz�H8V�K:.��G$��x�?�����/����M]@)��ֈ���ԝ�`cL�۳Bg���q�Մ�2d��%Sć)0dW�����A�N6�xB��C��z�Z���#���>���$�ڬ`�~�ܱ��S}i�qz� ���c���󩕬)gH�]�xN?���%���d��1I X{$~#�_r3��S��/�����%�k���΁��jMu~��j��^�Kƒ��a�ʶ���Z��7�qW���%
�����J���`l7h��ȓ��ꨣE�T4lk�A(��B��Aכ[&9 *}���G�lMwSɡ�ԫ��v@Z���Q��P%��]o(���
��5���ˊ.����3�gި~���F��%�E�W�J ��������B� �{��6�֎1@$�Hy�!��s�oj%]dQ
�/����|��s�!���T����(?(1h-�ݪ�k}aR�'��Br���}�Ɖx���a�>O��Pߗi��}�+��h�Gk�h�fr�P/���9/r"9��������bD��|y�Q0�`��8��ms�〉.��#��b�)�f�O@� �|�Ou}_�LȾ�}$(���6ՕOda�?6wP�W_�b:�R�iP�!�i^W�{?a������[%ϲ:h�(B�^"��X�����Ո����-UNn���p��,z����k|�����[�M+l�O��B��
%�<9<�+ˆ7HU�}�1"z��
�w[GN��Źpo-׹�s�J~����'[���+�����^.�N����H|�=�wy{����z�];o���u3x�Ԙ��D�z2$��`�H=�-!�WE��|"�a���͹~,��8Zd�\f�eHYūg�)=:�2�l�K�~� >�6��,@Dm9��� �iЁA��f,�t�=�Iy�!J��6w�xt8k;������vu��~�����\|�k�]�9�gjn;���z},��u�~�9a��R ���.���Q Mӳ�a�G{��$vQL�36�tYlS��F����"����F��7��ԗ��R����>M
��jWc�F�Hi&7< �<:�Ke�xI"�F��[FU��>;P���ٿ�@KΆ����2jtl.�D=W��D��uN�D��"h�ɯ̡8�4�u"������8ڸu�L	 �[����D�x�6����	�7�>��2���<kYt
 ULZ�5\����6�o��rh��ŀXA7ɞ� `�V�/��f��y��!k6�lE� [w�"&3g*g���`6�l�\	��ɼ���6��ZE���:�L��o[�Y-���ʱ�Sǚ+yk} �{)]�� �g��ڞ�9� ��m����Y���uՏ��"��]ӝ�6�r�F�*O~y�����(��գ����� .d������m����ڥ n� �Az�D��tC�MQ���B�~�eY]�D���Qp����@d�<J��ET�{��t��+�H%�lQ��'����e���=�L�QcV�U<`
Ш�J=b��?���-��-E:�?󬫥R�7�"�F�Z��o�;.S�z��7ó�P(ѻ����a�E�x�N�����L�(�Q���l���Kb�9��8�.ѝ0��a���*{4c���F�f��u���N�O�t.��Y���t�����ޫNg�l󺔨����p�F<ZWp߸n�b�#L��a�kƾ��#��pش�1�v�-߁B.(�Q�syzr��'ɢ�W��~]H!@/�:tGC�L��=�>%8e�5��p��h�ɦ*���p�D|HX�U������X�^�#+X@�y�S�ݰǂlP~YE��e{�'����7�n�|���zچ<�ێ��i������N8ʺY�<�]��/p��\�!h�Yx�E��I}d�A|���f��=�)�(�<�im_Н���2=��U@7;	d/��*KCe�5[�d�V�U4;�pL�WO%�� ����M�q
�O���τ�lF�mH��G/���z�:����Z=Qa�Ϸ5�L�CK�ڲ�3A$�L�$�%�Z�^�nRZ+s���u��6�a�\~��5'rFk�#�-��>��&�����#N���?�Ě�Y_w_~?�c :c��D-Z:��@R�H��46S�2��sv� ���ve�(M?�@���3��M��AM�뾳����D��̈́�p� �&j]�$E�=��>���n`����$J+8���Gh��ZÞ[��߷/�ǈ�~��`�<M�'";d��v�K�O��S3U"jg�s�{E�}T$�h~�0e'�6<p|����߰n��\�iu��&��HQJg�����}��F���˪Ӳ��"�	��2�$�2�Q�I-��,�|�Wag7�oB�Tg�ù����k���qT5�H�itmD�4���6^�h�s���v��9S����1��:zr�x�k���i��5���ܗ/ﳁ��-���k�P\�է�h�ʳZ~����F�.��p&4"n#C г陀i�R���6���6��3��m�|:��]��e�!t�L9�h��ſ�����o��Oulw�x����M�7vUI��iPK���6���<��R.�%m6$d��j���v������7��1��=kG�C�O͔\�&��!�	h�'q[���`z_@���6�)43�Q3�Y�Kø[c��蝸��u�=��ӻ)'���$��-�Z,�PG��w>��tڂ�'�|d溺y�g�tw4�AZ�P#� �e�H�N,`�7����S�b�E���Uk�Q�\��?���/r3��ֲ^U����y#��K���]n��[�����a�Ί�N�߱.&�04���j�6!���X$�=!C76y��}͛kl��ZRp��`�%C�%��E~�gw�O(�>*��i=m��T�>��v����ޣ����Cl�D�I�9-M��a�pu��#@IiP��z!��`��.>̽���^���ñk�	�B��늃MCj䟢�X�X�j��6@D�����Ky���
�Q̦��u��U�{��mΚY�@3���S�0'4Y��*��dR��L�c-��d�3X R�q��\M!w��L�����G%�-�ףuVW�8��UVS���?�$/䪲Ђ�Q�>sdk�{+wAg>�t��@�)��|-$p��8��f���̮�ӌ,�[��S�'�_"*�1�v���,:.���V)( 8���u&s��m�zbs㌁\�&�T/%� KN���&��Joپ��?���N�S2����5ƻT�o�D�! )��d'�[Q00�ֻ���M����Ŀ'O��t�e
�^2x�gfl#�N��1��i�=9��[�3�*W�؀]	`+��u3�0l)jΌ�&��U������+I��3kj��s����3����E�I+)&��ݬp�K�]_��A�Enf�=��'ՌS/I����s8�g�-F�&�:�r*}/��;��#��k���	`ɣװ��qR�漟߿��~�F\L֪br�Bi��t���Z
���� ��(��a/Q��J��e&��z��\���-�d�ͺ����&,`x{/
�k�����a�JaI��`f]�%��6by�l��uR'x��$(潉s���@�o���N1��<��Ay�u�M4<�p�wȋ����M������f�6x���*�1~q�ǘ���� p��p���	��@��.���;�?���ud�DJ���I�B���|�>��3�藀V����H��kX݊i3b��L�z���� ��Rє \�y�a��.|E�HF+>�e�YT��?P�芉(9��b�^Ѹ��W#+��oH>qCEod��]�&K�Ȕ�B�,6Q� R��d8��%�4��4� T o����3�_��PV����Mmʰ��!�z2�[��~��qᦈ!���NsOl��P�?��A�^��M4�L�
�J
�G����~�ˤ�����]u��2űw ���ֺ��O�p논���EjWd¦�^p%��q�J���7����,8�/�m9ԧ@���SU�3%o8�Di�Hۛ����l�yV1��A����e�a��%dr��k���'}�a��CiѢ|W�q���A�2�����t���[Hȟ(4,N�_�O���"��߰�눃xU'5���U�¾;��Biipƒ�<�e�!h�{��� f:9�YQ޾?�TX�K�ǝ;��w<�ڷ% �Q�1�o�2�rVj6Y�X�.d���b���:���#�Ąb���h�%�L�0fD:WN�+<I"�7��$e-})��fvSȝ�/^ ��؃��Ud#���uox�Ք�2���6�0�ٲ5�̽<���y��n�.�3��,�|��n��>M�u���;��9q�N[�G�W��@�ͯ�6/9�tWϢ����=y�9�>A��P�Q�f4ϣ���h�c�8bD��m�Y7�|��h��g�i��?Em]Ǯ�o%���qN�Cz��5�������d�ȴ����ŉ.%��Lr�?�g
y(�&�X{������1����:���l���NG��~���Hgt^b��=,����Cg@��M͝�����e�g������t�\��,c>'[���?t�*8�]�D�HM�MGqTw�_�(��r���z��u+�q��)�|��?�g"p�K��0r5�!դ����um�mÅ��@��h(*��(������+\)�Ԙvɡ{����^'��{�t��}�}���\ַ`5_�=ԛ^������w@)�
'2x��6�[+"�Z@���{����ky�ܔ�Խ��b zۘ��G��ʥ�ljH6�ن~���1���M5�����&^�a�I,p<���I���?"����l���8;K�I������Э��	H�e���ʰ?e%�g���֋V��Τ�lu}��H�`P�"�SP=B�<Pa����?����BܐO��qa���V�I%i�v��4p��Kr�^<����f��x'��	���p�lM���49�Tz�|*��pƓ��\�H���0꫑�2��+(6�f���L\�'Q�f��:���|(�g}�L�����tLO�����E�ז�8�j�5�o谐�;�{�����>1��n0�X��9�c-���{�C�5>����\ �[Z�u��4�7;=y���~�ϡ@��<XjZ���J�/�BG��Ӻ#e�@�W��/��w�fsI�Ef�!�6~ ��j�.��QHt��ak�A6w�~ ��lR_Z2�n�08�	OR$���O��a/��f�|�./'���y�1b�X5�T��x�ڒ��#9�#���7Z-E�@�J�6�ܭjJ�N=I���G�n��$�~�m���˔���+\���*̊�8r���^�V�]�G�6uط����jInˊ�A�g,��5���a���1�{T-�LnI�/$�D�gV���Z׹oƂf�1���2���Z�h�j����YJW���]�.��ʆwv�UCT ��/���ҶL}�!��y'x�Z
��G�"W�Ҩ���=��E�a=eg��f�b��X*��qF�R�8<���+��paT�7mB��7�ҭ���=l�Z� ��}#����S�'l!�5�Nj�[5E���Ѭq�1X�i�lJi�{wo���H���z���r	�
���c��3pEy��8	�:��EĒ�(���_s��e5�9!�6<5��~B6�0��d�A�OW��Dv3g����⁰*��4#GO5)Cz���b�v��I�-"P�6{ ����z��Fb�/��>�/�E�����x3�n�,��df)ĕ(L��
@�=HE=��wL��,=�=C���6R$�+uDFo���a�������u\;1���6_f�`5�	�.��g��n��#������w��������y����@$#G��y��'rD���g���k��D��,�%?�G���Rzd7��K����<Ui������
r�u�4V�S cծ{�����=ѩNS���x$�KI����\nU��ji���(���eO#ym	o!6�#�D�-E��~)���Z�`�>kZ��|G!�  �DӍ�߀��>]́�I���и�2�V8>1c�3N�x�	���rMCƾC�8�r�aD�G=�x������{��(��c2�3�>^1S�x)��߂ŋX)$t1
�!���Ҝ�n��:�AQh|y��O�g��wZ��,^!�@EA���;������JI@��nש�p�y	��|[���v���>,oWLd�3�jT@��%aJ�P*9�Xp��_������k��Yg�Ԋ�d6�F�S��]�,=yK�K)(x���2�`x�N�LB/��^D_���<�X���y,{�o[���$䨨'7�z��U�FNI	�ى��!�* '<ʦ����qW)��h�x� \Z�/H�SoS4&\�?љJ�2n�x3�g�G׽�-���S���� \Q��Gh)N\Z*��Yp��L�M��ȒJ���6��j�:A.�)�ga|Jb�.قU��գ���&e�g���r<!j��Έ_�l@��yU�V�{R�d�%����W.Ћ5*Ux�E|�h��MWy|����R��_^�`�]�FPӁ��m&~�	H`������z�l�397i��D@��iX������tg����#9Y��Q9�ߑ�uuw�`�-.�_���gc�~�5��a1���ۜwv�v���L�b�x��f������7��2��jQ�m�#��O�B��|q@#�Dzr��js�Xs���FaD�*t��@7*WS��?m��`@�0�U.Pf��i	���<�e�侓(���/����I9؆� �V�9�&?	X�Ү?y�bV4�����8V�J�G�l�g`�N�[���qI8��EgZ'6�6����A|"L���7 �wz�+����\�j�"���*�[N4b��O�/��������Խ����v��?�������~j�W���#�BbuX7T�+��{T�?M�A'\w'1��� �D�⥢�԰0�c�ya���#�Ɏ��|�&��x�3w nLtdQ��_%ƒ{��c!3:W���׫�[�£�LtQ�IUVV���A��##�+��G!R���l�؃GH�0�1�UH\�X��Mrt ��<�$�A�I�ܿ�������8G�dj���
ސ|��࿈������$�_2.�B�����)q5��s�"n�T��|�U�8Oޘ�ׇkC��I�,fz��g��b���'\!h��5���b��I���$N~���n���y���"2��F{�&>�_�9.��&&�Be?�,�����mG�c� �Fa��xgH��#Ib���(F�����f��c!YEW�����"��T��qI��z�~�"�������̻0.`�H�/=1_�z-0We�ā����j��q��J-͢;��٨:l9�C�L}b�n�k=�� 3�����V~�j���L����wӀ#io�Z����Y��/C���Q�/�,_����^M�6�N�������l�|;a�1K;���؅P?	l�w�������f�5`�����	�
sF���d�lĲv���lj=ʵ���)o��I��k��_�/�'a)��$-K�_��u�9t�(.�hf�/�@vg�O�6�8�i5�B{�"��e��Z\�J�i��*�x�W��kݤ���������*BƔ�65҆�v�%
$��̷{Zt�9\Sc~Jw���g�P�+�;������gmp�z�5�s��?���W��)��"=U@���#S$�9K�X'���>F�`�.F���$Ld��ԂU��&(ㄤz��J^9�~���N�v�3�:��7�j'�Ы��]k����M+�;�B��s��e�f�W� ��v�����ٓ�5�2� Dj�qx5�\*��m$֙[�t�s�3�2�*�pO=�bFL�n *m4��EӀd�N��aL������(L��`M��}P�8������� ���W��Pt�ӻcg�,��D�����Q)ݶkE�q�J,a��I��-!�7�������@0�(M�e���aídz�?�^쁡�i:�g!����,aq����K]��UuیC�BP�;�h�?_����_�z�/{�(���$Y��1R���Ih�_fWr�&}j��L J�F���:K�^�m�w�QC��pN�kFe���E~
=��|�����sH�X��ܵ�E��&gG��iҵ'w9hl��Q��Hބ�Qw��M���b�Z��Uh���>�5�_�ċT��	B�Ս"�~d�3�=}����sf:E?���#��Њ5�'m6���0�Sô�p�d�V�����d�=ܝ(f<(��R�I�=yp����;��<gN#Tu$:t�_�Gc�|f�AєY�8�&�	�0
c	ۗ]0J����T��
j3Ķ�u����-�b{��ة��ۖ���ݾ�Җ��Vz�5~�-K_�!׬�����V�����v�:�Xz$��$tPϧ+ekv	7��yaI����d�<��W���EQz���=��r&�S�G]����V;���y�$�q("�����Y0�6��S��yb�`����r8/��8U���1lo;y޹�Wғ]�<h7�%�e�����{Lƭ�Mo�/���U�@څ�ᄿ�yL*���F!��_O {2i �HпKq���O<ݥ1� �m Z(tO�k/U{-�}d��~{>8�-TN;��N臻���a�I�B,�����p��y{`� t��W�<��/c�9�^���;�7}^v&S��qI ��J�V��:��i ���e:�Pn��}p䕲uYMO�]j�3��Hk���o��0��Q��M7��"9����iNX���~��%(E��[9a5���ZF'���9���e"�a��1�@'�_��Om�Ol(���^iM��f5I�W�؛r�.�<�STI����SB|k�(�Uc<��6�3�^A�_.x���˹8Q��Uq��ӱN��mꝖV-���a!$kVs?&D��R3���鬮�q�qm�[]<��6	b0`Ys��s��� �Cٱ��-�C.�:5��~�m��P���ɝ;���{�/�0rj�:JYNY9�k@�Z+z7�@��fJޚT��R4�9�<�>����I���_�Z��ɚ3�&Ne���J}w�~�����<{^_�ȳY���� �y�9L֥M�)�֐�9�����f���/X�
u��ԉ�u�p(��*C ���e�ucY̶�|�����a��C�n��� 4����v�Q�F��7�5BH������i
uVc8��{?��\�n��k������H�Z/��	��e:^��u�B����
���S%p����dS��{h��()W�=�
zE���G_U�rGm��TdS�>N���0�������&��|��&�8�@S��=��Z��E�m�h��[^���T��A��
As^ 4];nk�Xܝw�M~���}�/`<@�����O���.mk/��!R�&��؈��MW���� qbMOظ�"2�DĈ�E�hXR�;�O�����u��`��^?pM�v����>��uD���l��;�� �����n�zz\�F�� Ų4p�%LyM��kҹh�T<�-�f��������fRө�G�ʅ�bș�i��&V��Zm5ߵ�`m�^)�M!�7����{����cb-�9���m����p���B`�T�d ?3�WhD�9�)��
������NF/���8����+HH$��f�5�01f�S1N��E�PU�M���N��֣�+��(K�,���۳Ѕ)@�S1��C�?�ͨ&��wK\�(΅rϢÂ���%��w�ƢX���2Jݾ�5t �+~�ZL,򓄲�C�L����V�f%J�h��;M^\^�<wW<ň���L��oKQ(D[�
��qеp�':�o,?��IA�%ם\!���5�K�p�qj��J�f(�[�6���ݱ��3~1v�/T��=A��[�5�E��1�Z�TKG��@�# ͺw���,���p#�Ƨj��P��Ly��_��w��T㼜�N7�o4�����	������6z��0��4CI�x"o�Ē��$g:�sZ��FWU�YJÂ�p3�9�p�����y�w����P}�/)W��<5y�?$��>��ZI�7jY��a�yO{6��Cj<lr��5>/��u�t�a����=� G$�I~?�z$kG�h!�J� ���� B��P�TQ�.�ɯ ���G��3����!����p!]A20^����O�eCx]�G�/	�{
��v�� �������#��z��|S����J�䍾g�)�pJx�1hʌ@�Q��9
�7�����Tf�{�A�z�|�@� �΄�ǟr!c�n��Y�#K�<J���w��c̸�����}����mXV�/��<@mp��΂T/ݢ���������t0]a/aU���QL��>rϱm��ޠ �6S�;�Z��F���()~>��m�(����"�D@Obh���ٕ=���9WaFvTWȶ�
7�1�|�M'C�Tq�uҠ~�A��k¾���������?f�Ԁ��Im`&�w�T�Sg�D�H��G�2���Ә-�>������|йӸP��a|:o���������,�
k�8A�ܥ*�ųOc�׉,V�n=�4����H�9��q���ر�~`�;�|��[�"�/�%���s�`V�t��­����t��Ʊ!>�;&L$�f76f��0�5���򕹓|���՗Rה��5g�\]��I�l���{��;
^o��^����Ya���nM�J��������Op{�bx�D'�4=ri�P1����J>�����ئB��f*�U�1��[d}���ҁ�!x�5�k*���>��ӄq��{$i�A����	�4)�
z"� R���!���'�T��#��#L�ɉ ~�(�q�n�XdD����~E�]�k��{���6���=��	wD�;	z�7��ӌ��_߱=uŎ�O>x�
��i����'�9hw�=ߌT�12uR��6�Vֆ�D�e�_r��'������ʊ�=}��wO>�r/σ�ڶ��|��;����.%ꤹGUc��������{'Q���v%-��RY(�k���VBh��}��7V����C@bB(����-bV��rU`s5c���FS[c�ԅ�V�����0���|N>{f�"]0cv�ED��7zzߠ�
;gDo�hܱ���PaU�t��>�(�T��3Bp�{;&�)~�C.v�$|��ݠ�]Wa�U�|!��6�g�����6B_�6�q��BTI�a�"�����/*���`9ò^s�m-�����V��/�OϮG�~@�U�5l(b$Y^�Ƴy�qV`
[��,`2������Y�۰���Sg@w��=�l�X��͠	��j:�do���{��<�����NvP�W��h��"�H~������Cy�Z�
+�wmy��8��E��Tj9-�J4*c}ǭO#}���b�%Z?Č�@�LӨH�I�F�fu��'�M���&�)���|Ϋ�~�%_�$��8��y�U}�;q��Ӡ�[k�Z�K�3���=j���oĪ�!�I���-x���"b��h<V���jv���H���6>9j�C�rx�����pY���r��~��z��ldD�I��}M�Ĕ�Bq���n"��7a��	G"��+n�=UdC��(���HDyn��}�k��ɣ\�J��^����C�*{��9����Qn�XXj	��8!�e'�%���=��g�}�_����ᗪuN+8N��}u�� _Zg����%�����,ܤA���[���o�K��
4���U�hyؙ&�]�Bɠ����~�=f3'cL<��A�Ʃ��ƠY
�k���oR��g�r{��â�]���2W&ծM���U�a�R���}dV�`%��~("��6+bE�ȹ�S�L����ޒn0��"(�/��B���y`�:�pt�+2�J" �ᆕ	jI|���Ź�e{�������=����y���j��Υ����w�#ΒbI��o0�X}th�2���&���'�o��� <�	3���>F?[�"�/��U=��e�&&�������J��1���D¯,s���gHmV&�7���٣��@��;	��ݕc7'S��A�*9+�����Ғ,�
��Z�������Xm���p�
V��28��#�Ơ����wyמfr3���{\?Na�ަBR-,g��*�����L߻褨����EBJ�d�������A؇�ʷ2<D��'��~��<�z�Z�L�Q}ɉh_ŉQI��Vu��_a�?x�x��S�%�}�iǒ�j������ ��G����+����4r!�޷�1h�a���'��d�Wޭzы8��;��T_�VMW�H�@g{�nϥ�,��shX��p��-����ˁ��>Lj ���M:���s�hqɻ�Pހl�j_���i�H5��BY���:�Zg���8��J�r6��X�]+�7�B��������d��u g��Xw�i�0il����.���:An�gU)V����։*lBP?�UW��*
0�S����%0�]��*����;&��^��U	$�^?6)�&�lc�7�G�h����Rw��[�o��+�R�c~u���G]�� ȝ���F��_��ߠ�nIc3u�n�\[G��M�Mw	�0��u�-��l�OKH��=��[
��m�<���i^E�� �+���̥��^��W��;	նlv��,��C�G�c�Ui����<����5�����b�����a�J�����`���]5�������?6�RiW�5.Gq�kӣ(�0.K��rO~��*�|j�����u�_i�$Z��G~\�`�p�=����
)�q/ޖa�#�aj\"Ŀ����Z3�L�||���>��g^��0o�q���E��.Z�⹛d�z�|���o`�:#�+����ڔlJ}��bR�4�p$����E���CQ�Q�Y,8AQ�f�6�[K	N�f�nL���EǦ;�o؞*\���'�ꬵ_����	`�7<~��ojt�%��4ߔ�
�~�ǖr)7��,�EPD��K�-2�j�5A�$� ��C?G@�P�OF�P�e�z�T��'0�a^����(���?�:���c��D�a���
�~7�l�DN�d���>G!/Nϧ`tCڶ���QϠwF��2>�[F|<������V�p��/R��+K�9�O�L��,�g6�
�OS,�B��x���G�����`�H��/�ǥ{��Z�J���)C�6(+�\h�#�|��.2��4xx�J�h�:�c�f�ؐ\]�ia�4@ޙ=:��I����<����߇�Ж�+*���~&w��y��2U�9���mT4v/9�³�����7����zz񌲆��KQgƭA�B`��{��*����ϰ#��m:�q��	`ŞV����#P9W�Y�O;Gӟ����	"�A'�^8v�����u��#�4U���4P����2��0�2�����\5��R� �O�fQ�t@d��TO3CZ2�fSO�KA�����K�jݸd�滒��r(����t�˭�h/� x���΄�}|���/��� �dKG���9��;0�o|�'� ^A��Aw]�}ҨsO��V�z#�����ջ���V
��3uM�����2J�����Ҙ��a�L��D6��B$����+��ܻIs9ם���@��1,j!�L�yG��s�˗�F����l�3��-��K>C�{���S@�s��4
����1���sE�	����;�%�I�Z�R8� 1n���h0s��2���6�b��;H���z�g۰.�������h
y�����I���)�ng�w�:JPRT"��������\xK�9��W����H��&��P����'=%8#G�~�r���D���ł1<��>�ˏE���#Q���EPJ���6���@�w�(0�?HSI�c��ȴ�yF�jADmw-��ĵ�������*�X�@��iY�6�J]����W:9�\����:=������U���M��i�˱�͸	j�YB�YY����y��JA?�]Z�����PpS�	��i�Dl-1���:��#l�
��t���~a��o��bq��V�MFP�T#�H&�x�-��3��HdςEIE�CC���9ge�Sezf���j�w�
�K�o�]�`�{24��a�怩�W7�j���]&6!�g��-�e�n��1;ݩzFN}�}ޕrw^-"]�h��_˸K��xӫ�EC����J�@����֌���,���pb��}�x��vG�^E��ޱߔ5���W]%0�D�N��
i/��;�>{u�x��+���"������-�%��	v�"X���l���W@qz#u1)���5�B��u��K�N�%?�S�a�Q����E����+�4� �F�̑B��gM&?B�������3��4Aͩ$����q�>h���P�ue�X�R�@SÑV�F���C)�G����~DȐᎬ���Uڐ�7�?+T�I5Dn��DL�� �U}�:�;�a9ɘhh0�ORu�T ���Ƹ�Ѳ��1�o��k*;�0o��a��������?�s�������è��GƆ�|��K��Z�;��!��8+Z
;�3�6�C5���{��\���;sp(��O�)�o�v>*~�ө*&�g�*�K�m��E)]�|'M��W�����*��R4~.M>��ʀ�:�Y;t�b!�[��Lims��,�Q�S8�t�
������mZb{�s�'�Z��*4N�qI'���KC����)�����-�0����am<�欓�:cϰT�6қn�<�]�����Q- ��)���`Ѣ��t�_a�<���~v�%w��)u����=��qL6�6��k?�r��>�l\ $�v��Y�0h\ %�o%#�Ajh�� �²dؒ����J[�Y��.�ޫY�����CN�� ���UIy՘�mM��ƔѨ��~p��v�D��x9���5��+Y�r��Œ։1E "�$��a~k�nF�E�O�-9i�Z9HV�K5��6��wڡ�^+�����0��*�ko*����AQœ�P�5u\B�q|���]M�~X���d��	S�P��p
����c:sr�d�$�ʬ�A���p�eJ�׌hd4����h5.��(+iA!�?Cc�ć8���T.�N���|���/9�
р�����j��~�ò���$�-��c�R�/TnE�ܶ�ˑ�c��83t&�}��l��
����md�B�
�HR�Y���&ģ���+����s����� p�.ڭ����r/�zڮِ����Zp��K��χ/Gk�d���|5�1�H/`���j�$�8߰�o��A�,
#�cV!��yF�щh˙�A�d���TM��~�zy� ����b�%vx����Qf�P��:�%	�X	��06ì���3ĝ�W�����ꥅ-� 98�ı7��6���pf������F
��0I->��G�x_?(Ƀ��Z��",8
�L/3u�/W�YI��LQea ���ܺ}��-�Ǥ�b�w���R���Q�<�����Eh��O��^+�M頾���B�~*d�� 5���]T�Xj�Mw%����]9���q�e���8�/��d2F�a;�vȢo�3<I#�-��cuڀV�O:
75m����t�=z�T2~��=Z�L/]Sw�u/x'T�70������"�:�n�z��acjKI)���������Qf-eYՀ�k�
<�5z�����R�>/r}��t���AX��x2��S/�A?AF�se\�iv��P{�����YK뱜�(ί����ژ�ś���pF�m�&C���nH�;�C	c<�٭!J=8���B��c0�?^asr1����<c����Sd:�C<�v�~�X ̷ �}�=��!���NpB��=c�ՙ�3�p��(��UVr������VңxVꥑ��N��հ�[��c�~Mb����d���4[!�m<�½A'a0ED�����tLa��q��@�	#�Tx�b�� �i�N�8�Iil�)NG���)Ю��H�@�N�m���ג|�~�m��� =s�4��m��D��l�A�����<d�1�6������z����������	CX�`=u��(i@ r����Wa��^E��Ym��*��@��-"Z���1��(��>aa�f�M�� 
Q;%�&V䉣�3��D�t,
��qTLד6�r�U�YK�\��St��~�||��N9x��9k���0+�ȳ��4�qN�l��tkE�����@Bо�1�cS����=+BB�krQ�l!:Y��/�'_`g,R �t�"hw8y�&o+�k��z�7��S�k��*�u�׳���u�K�>�c��=,�!��b�ۡtY[�w��N��qNp?���~9mhDZ:+�+U�=�fwc"�iڮWpb�_Fǹ�	]U�;�i�8�2�5}1��l`��������& `&��I��A�����{��H�ʆ�����L;�-�[s��� x޿�$Qڤ)�ߒ�WF�����R�8��D�0�^��J<ZÛ���	|E1��n�l�5��c�H�ދP��i(�0N�(�w���q"�
�Ϻ��I�������1K��#����^�{���NU�� ��}�0����y�Jʼ�S�}�;�M�5؆;����6BtulBD"(�[�b4���ɤB�$�FĎC��s/�q�����x'��
�x�*j��Do�~�Ѯ{h�Ws�~f����HM~�ܵE��fЌ����yFK m�v����NuY;ڮ9���Lb  P7l�LbX���@�#���v�Wb$˃�Cx�R���)�J���O1c��H~(�
g�Cn,f���Ucv�&<��k�ꐔ�z��g�bF�u�ėm]E�ƹw�q�ӭ�����D��oɢ�G�q���7M�֎��(uM*�K�5`�����wk?f��PBs@ɉ��N��v)�݌�P�����v^��݌v���F�r�Ũ���䁎�,��oDl�4� �M�aGI��L�}Eq{0U��I�n�YT=�IQ��?��:H���& ����E�} ӡ�ȇ�zbgVV��x��L�P��B�
԰��E��s��H���C�����[��c1�. 0�����x�p�v��� m��M�� ��J 
�o�qt��u�����j������"B6��lD:`���+�7o�k=2��YTF|�X3��T�S�h���\�`[���8~ז��hx� »��PN��nU �9���4uYE��m�}����^�R`����dxA�vЖ#� M�����``�@�;k.���:����"���|;��s�ޫ*�tUࣗf6M���&V �*��:Ցj5E:�C�gƘ�@o�
��Ϊ�F9B��G���AK��P�y���_��Z�q!���9�}j�F�^|��[��	S�2u��-w?~O�e���O���h)J���!����r���c4ReW�x�^���^w�F�7�lC6m҇�jY/�L~��=��G��@�h4I�+���a�|d��E�!�eQ�w]w$c�.&�n�Y3 Ә I;\(}h5���YN�on�H?�����h�ңʢO��a���Ө��v"
���ׂDpr�!��L6xԂ�&��	#�w�5h���v����N[Ѳ�)�+j0�ϗ�6qg��ʴ�3
+*`���DR�4@�O��X�F�Rr�2qčw�<n���gq��&�a��pf�	�<�[�(�"���g�!� �4)�дm��}'�<R�A�AQA!7Gf�TJ7R�-e%A�r}��1����W8%�O�����j����/*n\�L���w��<�-��~�Նv���M����e��;xܣ$����vu#bV��}�U.�g���fML
������?��quo�<Or,;�i���$�bwI;�DQpH*zM�-gTƭ�g^&l�1���(�ȿ#���0��2<<��lƸ��_N�d��H��E��NAM�_mU�歧�-v�n�n�h���`A���+j���]���I��:�*���!��=���|�{��<��M�X* Dj3��fI��(�>>���ɀ��T�^
�薨�5.��
�(�������&-#���!:	�y¿��SoZ$J̢�w�7ITI�D�y���5ؾ�Un��0��|M�S˶\{��:}�)��mIo�p������_��-�ӭ��~�b흺,�bgԽ��
�˰�7XC�ԝ0�ɚ�b�͜�X�+�}u�+�.EiBQ�@g���r���� �,��{oƠ��|����ϩd�k�7eJ[�����GYI�>Pc{ܰ���]������e��Z�4t���ի���-���/ñ��8j(ň��P�����Æ=q?H�K�pu�s�Փ�[A��x��AH��\��{E�p�^@���@�4LRy�$D�]v��A��#�C��oE��w����9�\/ܴp!qA*s]����5@�����'�#~���[R`�ɡ��=ъf��d]�l&�e2���t(��i����nɴ�:u� �C�J�|����X��+eo�%!O�����n�P�yS���1�Pz��:�|',v-_RS�ũ�}EE����O�!���|�8O��1����87���s��AI������/�[XA�H)�F�رF��7�#އ�gl9?0⛰�߭�0�.ַ �Ԫ'U���ƾc�� �}�'�!�)^��R������jA�� ����N-'+oC�jZpf���o�ؓ��I�q�:��n$�a�67XQ�.0�.��C������ Z��9¼Ȭd��Y��R��xUelƒ�O��������,K���,N$��u:�5��_���s�M�0�t��Cz�x�.:Ś��Hn}���(�I��56�\�W��.A+E��F�� �vD�m��H"t ��Ե�ɒA_.-�8Rb���x1JT��q0��p����[g��tmjx�2��
�4�%q���˙C�W_� �h�u&��I�*^�Qd)�ϖC�"��΃؝��!R��$��q/Q�I�~���u,[���Ŭ�' ��XQ���c&(�*���"����6-��V�;�l��>���i��A��"A�����R�{}�������P�z�����}��1���/��z��N�l�V���c��ZJ�����A�ƣF��g%��Gb6��u�E	��'v����sّ5$'r���6J�чe'{Μs@��Ж��|>����w-�����
�k2>����� �fșq�X��ȱ,<�;�0��	r�N�Zq-K'�H�z���r��[U��2�^jsS����&��q�����c�MV�U�l�o�����>�������
?�PI��aĨ�*�c�m�<��ө�|�9�3!�;Jk��y��
PtB[�ģ���2A��N�ŉ�V�{f`�M��F(�Q�o���tSo0���<\�M�6|t�� ���à�Y�eD�~�ɇ�q���51Hi�ZP�Z�'�%�j��`���y�5�C�Z�癴�����-S��+�u3/�&RPߏ��M�fu�*�f-�xL	0�/�p�ϲ��
��kH���cC�N4���F�2��A�nxk~���W('��(>jSy�&E:��3�#ݔ�\��dn��5	�̺#`�w���E����4����c�|��[]��e�:�) =� L:����?|2����<V��	�kF�f�5�p����v�z48D�"'п'*1��p����ĖM��a��rڥq_L5p���7qZ���'��B�����\�KC��:�ν�n��Z�|�K���^<�!mD��MWe�w�e��(�a_�5�P��T��SY��8� �!�-���B�[H����b>���:����/!B���{��@�@����o��9C�V]gZsFb�}�Q_��,� �)���m���3]Åa0��U�W	����]k�$斱[���5�� C� Q�;����7,c���Q)�*�YVl���6�}���v�g�6"PV��Z�z����Հ�W3��!�A��<(��Y���6o�� w�[���y�[h�(�+�O/�
���*8���%�BH���t�L�9�d^��n_�u���gO��:w��~��hYl�I�QQ�-���dTS���\(֬h=Sl ��{o7�4�*ї�{��Z��T�� )�/ a�2�B|��
>9�L`/���1� gc=X:����z�6���D�p��7
$ų�t���͵ڴ����zR�U�	5�N��H�]J'o���#�����C��#������Je�v0�A���gK�7�����r^BQJV��V��ѧ��M�>}�eK������RV5��V6�� ,Qp�F0�2���+��v.�u鵹��� ��2~HG���`�l	Bz� �����1B������s�:+��-#V������{�ֱ|rY�L�^���0>�z��B>Fl"�.��׬��Q{�u��A�-��kY|0�9�H��^�z=�.�c����CF��h����hO�X�r���������_��f�"��?y��Z����7�CZ��y��t.fbu#O��x��-�L�z��f�OM�V2��	K�а@W�QV0�eu��˕^R]�C3Уj��k�4V&���x,f6��]���V�ߚzdN쨭�|�:��$ͥ�SLڵ"�͉i����z���(��v��V�M�b���� ��vA��7��z�[ ��P�ri���
���~X��QO�������6X�iZYa;@�/9�S5'�fz4b6�U�Y��3��P��4�}6�`��$��ZK�}P�5i�w%݊|4>�(o7J9p�/�^�'U�U�
Y�-�+nZe�@�ٍ�`�|WaW75�㏆c�soPpy�є����_eV��%"Z�m\�Ӷh�ʙĪ���H0{�a�v��)���I�N
�� ����}��LQ�~�0pe�J��ן"��y1��)� 槦K�Z�̖�g�ȵ���-�S�=otzF��D��ܱ6
p��l��I(D�40z�����R��U��e�u����T�jo,�ޟ��&{�'��0�����Y%����c�ѓ\"{�ܣ�i`�ޘ�
6k�u�᩵��lR�$�PF2Af�o�r�1��i�t�D4��af<m��v��D�-Qȅ��f�>l�ܪ��U+K�e�0A����I_��.&�O�e�r�$�.Ƚ�y��.UoF�\�����Z�c��+����dq�'�L�e��E�2�H����6�q�	c�D�B�����!���3_�.�u��J������ui��c^��9v b���!�5P �\��^��Y��jCD� RX�Z�K���ɛn���,��7��{MV�B�����#:qGɎ�ڏ҈�5"�%�{��{�L�����K&�E��}���
��t�	$����i�^ψ����6�}?��2��S�j쀐U�1����)�H�����P��;-� M��2p�H&��9w��̵��Y��y�ҝ֗%uûf')3KcA�v��I�D�ע>�RJ?���я�������a
y�7�wo3��K�*#���?V��A���ꍋ�J^W�NA#p��5�;!BO�W�� G�i(�N9�7٫���Üfٖ�����V�B|���O�T��8�Nc�~Vc�Z-Ѭ�ȡ	����V5ǵ�H�>�N�,(ەxy�h1�e��k5�&��\�G�ØY��u�R��f4M��8���� _����r���>�ՃD��M4�� Z�#+�rR �-�;���~�0��n$Pf� ��(��Xf+f+6���i�%�5���A������D�x�����h�L}�"ȼ&ve��R���澦�U0 <A�`�Ȧ+�v�B�1@�q=Y�fl޾3��Ʌ�ܟ�W�H�2`Gȇ�<]��E'�ذp�l��8�v4S�����:f{LW0w����mY�V�#|�;J��w�PX����A�� ��u�����y*Pwi��O����9Nɧ����Ǎ�#.��e�{3O(3Fx,�#�=)�b8��_��_������ٜN�n���3p�Q�/�$�z�t[�uw�۫�g��kU��h���J�K�D�+�� Nd�:�x/�DG�m���PY��E�|}��c�S��G.��M��]{�F�����:{���M�Z{ȴ�\����*o,��K�n�e�#����p��_����r# �f�Q���Fvec���b�}���N�Y� Z{h5*6QcC���B�i����r���X�����hvH��$�N�XȖ��}H�4;x��Jk��m�Џls���e�Ġ�)�����J��`̔0O	�
��7�Z��M���RdX�{�T�n�9O�%(�>2m�Q\��"x���`�3�b��	�U��ϳ⣽�s_�����'/ ��dɾ]j����eW.��v����'I�v-�a4mDz�!jx�o��ɇ[j�#A�۸�Z�s;1 ���� 2����ZJ�_�g�h����_�	FK�qd��FZ`�"yt}����×a�)i ���ẙ8O�#��r����r�F��=�R�\��s4Px�B��P�$��6�'�v�.� �꣗���ے�1�����!ǒ�m��w�v�96���b������N�5wS�L�T��#�����7��!�q�BC<�ɲ
�텝M���}���x��꥟�;~e�	ΥM1�s֖�ͬA��.�w
B/�����x�orUa�}K3�/2ܵ18�\���5�9QXiC������<%��~�!"�3���i�}�B��i��veY��}�Z�٦��>�z!���ʈ�m,�BoSn��||��b��Cu���c6�ZB��NQH1���@�q�V��@D͜�����>VZ��t>���^q�V�8�FɨL���U�O�����_δ��ڎ���0V"�>��(-Wp�Q UW��hᨐ�F��GB�?�ϴy�Ɂ�_���f��x�_c��b��쫫��j�]�=o����i��[=������W<GѬ꺧ݟ��6��j%�Ҙ�K?� 2��jm�Nn��;Cx{޷B�n�KXk���z>l��}uK����4#_.�D⮑��ё�|Xm�_�C01`d0L�;����/#ڿ� d+xq]�}�+X��%�^���ۼn��O%ݒ�<����9W�A{_V��y)�W�^�,��Nt;<B]��u_g�Aj���5D�\�~ٝ��@�:���^�'��h�_;��-�������m��/�[�DWJ�l��|d�?��x�xf���и9(�ī�!ijw����V�����H`fo��󨊛~�$`ZC2R��٢>�j�k'wڃ�*�c�4�m��=��H�_���Zg��_f;��"�m�Y8��#�x~zL�����FmOq�җ�c�V#t���\��eE,�HA�q��
NS���O��5LEh��G����frߛg�<U��ϗ�0�-�^��r�Y)�Jv��/���Ĉ��Y�^o8�s�]�%`VU}���bNtfH��T��A��6�����kp`���U�,�����B�+k������w,7�1;�_{���4���_G5��>�0T�e�(�[F�xʣ��C�'����h�Q�Y��Q���OŉR��@�9K���-=��A%X�eӲ/^!,z��s*�ˉ�~��	�,��k>�n�>�Q�d�4���T�0m9�*�a������_"ũq�	�Zc�`��Ȣ�}9�	�gM6��h�d�����{	�ʆ�j�*�k���q)D�U�+�J��o��߈1��BO�	U�n�^%�D�O���8��w`���un7s�X���6��@~
P��g��W���m��������[���D�u6v�l�g.����d_�f�9�Y�(v#�(��?\�w�k�n:'��E��<&t���@y��z�~sE\�\@��A�̋ν6 �-�}Ak�BA7Rҵ�b�1�lͻ�V�؛&{�x�X��i���HD��̝Cl�Jv�/�J/�l���˳�~`�����V+��M{U2���P�r�y�f�E[ی�&3k*�r�O�s����u8t���mB���}�z���ZH��w�l6ې�h&
�H�-�d��VRqvb�u(�����
������rrkb�nJt�;��M�{�~c �t��	܉����wq>hJ�_�;��'F7��8)>����jr����X�����:�ח����qA�0�ʄ�X�n)��<��F��޾q���G�3�Y�����pj�5�b����/���O�L��~�R���L`�c:�� V-6X	vu��3����l}D�ٞd�+j�m��cz�fǯ�������Y�RЎ�L[wtm��,QO[+t����͝�̞q���/Q�˕Z����>��ܞo:���.� ,2�NE6��Ƀls���<n}�5�پ��P6�e���1�R�9mr\�� �s�Y���1@��L����M������u]�ET���e���h2�4C�3 �N#� D�w���x�l��L�)0��R����yAm�ף1�hQ�
;b���6�񯃇�۲e�Z}EO�a�J�.�v˒���x�X�}���y����dj���G�.ZB��@�b#D[�՞����<��`���[q%�zb;�q����7��"��b��9W�ˤ>��Lq]�� ��8C�8�LǼ��&���q�4}:g����H��~�A+6:S�;.<^��U����O�i|���.�`�l�]���I{����ޔg�p�a�{~q3_�A�z �b�t�β��Vh�@��gO��st<ܑ�������{[=��ܧ��뢲�R5�Q���W�;�>tqG�l�"s�-��Z�ev�D�(���Ya�r�i��L��,s����/��*�r��,fs����++�1s�ņ��W�4�!+���&�z�g���PGCv2���"[.�����dt8C_G�cUz�N��b�mC�v���c��^�Y�!~��$9A�1+��ҫ�ǠH��'�:Bf����>1�!?�W�M1�7��m=���̬�[� M��#��J��T�R��m����_�c��础Рu�M�X�KЋ`�ۂh���%BⵡB����0j�nLmC�]�n�Z>Ɲ{{���u	#Z���ѿ���xs�L��K�Tc�\z��IN\˨�0�gh��V3�Z� �+%~��h���BӤ�웚q�Ҏ�"��lF�t���窟�I3�EMx��b�됪9?T��Ե�t\m�� $d&	<^uT�ܑ~�Ũ͓Њ�áE������>V�^P�0E={���C�P#l��S֐������z����sǗ���5�xs̊�����v�r,0;%V[=�t디U��?�SԶ�b~�0�'�U;���['�Dr���)QOm<����}��"�PE�"K�r�5G,������Rd�:%6�X�Q���Pı��dRtcrP����K��N4�ne� ��ϕs��ˍ��ࡎ7��3}M�"��V���<���>���P���`%RwG�(V���3�ݡ��� �[0��_��Stl�1��d�5�3�3H\�d��f�6���핌�Ņ���,�N�#�M��>�����j>'�q���w��N�2�v����P�I��3�N���&++�VIm7�(5Py�������-ն�l��b����f��" ��ں��|u�ݰ�k͌���F 	���9@OE��I��E7v0����e
��՗�;�G53p�^7T'e����x��D�� |֝4-��Y�An]6��3�(��(�u�lM���AD��}�����R� 7�f�d�T��z�����%�Jd;��E���@��|��$#%ۅ�Pky�Zo��X-��_�����:������|K\�+�
8u^�:A)I��'�r��'��U���t�m�-�����~���0Z�Σ)�!�D(�M����8�{�:��Zqf�2Z�eZ�h9{;VZZ�:	�`U���tn/�����

�w�e�;�VY#�'�$G�h���;[���NΞ�c�ڼb�329?�sb�Z	�	�~f�2���yƋ�w�c�\r_LMT[�y���%��R��7��c��<��8U�ĽЧ����u�f�x �$+t�e�Β�����S���p:��0e�i�H�����_r-$S�;�V�x�^Wj,${�D�o����aJ�3����,���Aw�23&�I-~�f��$$E���§I70֨�Y;ث�4KjL@L�� �� `I�E@
W2�"cQ2MR����j3M�m�,�b�np�e���1M��aDI��Y� �k"�y���O��,�?5X��!�MY���0��OO�^M_ƣ�=���P����T���V�z�z�?� �*��w@--A��>D�jU�'d�ӟ"����v� �o��?���S�N�+ٙ?�(O�!vgE��;X���O0�_c`�m@#�s1'��K
�E^�&���Me3�3�Ym��%��&-m]���Zi�C����`S-�S�A�4�Ku�^@��y�w5�0+3�@]����/��ǩ��Ȁ4Zu�/�W.�I�P�b��b��:?H���������?���S5^.��YE�0뇩/��r�Z�U��'�Y��<��{t�ơZ��TQ,��@#G�|���-y����r����C�%��
>0��������vY�Z�e�
�1x��b͘��0�?�I��4�����'�A �����UM)��wXG�o�8_�R�Ҡ�	{���fJt��Zf��������JD$o��<i����.s�[	�>������nN�@L�w�t����l{����+t3�S�<������0��%Ri��r�Zd������!�l�d�������g2?���0�����@��M[j����	��e��k�ࢽ�\�H	WU9=Z�@��.D��Mʖ �(MO���^n�tZ�𹠷�I�3�\�u�����n���<p]�
���������] h�Ym����E��g�|�|��+�q�AY�L�J^���a�ݣ�^M�e&7殷ݢt1f�k�2���{�S������L�ܿ�K�������V�?����O�H���O��k�,�%���r@��0�Z*e,jp�=��э z\��؄*2�VAY~����Z��0�e4/��
g�R��ʾMZ|x8u?U�P_�(���9�LI��󶳣�,:�GpM����u�0�'�T�fjPx�*'�9@�ĿH��f����ua��uR��g��jw+}�Ǯ�.nSW���|	~�a<BW:�#�	.#	��Z'��%+~k�B�S�B�$4� �K͋|Յ�&
�?����0�\E�զN��3Ƨ�����e��.�Yk|��$�������hQ���*$��lȒ͢�$���������χH��֣p��������5��w?D�h�@����Ʃ�ڳ�oǟD03��S���O(���tj��b���6�\�A��j���ӎD��2��,ҏ���i=-_xڢ{vʿ�� f�!��2E_�!�~׆��X޴�b�I����Uv��<@U:�����QM����i���Ocp�<���.��,�0nB�@��9=E���>6	�`��i0��\����L����k��:�����!��)�W=��©�W#3�Q��_�(CD�Bg���A�������>n��A��,u�����h��tp���X߇�F1[_[&�"����$O����g���_՛��k�/*��i��	�Ϟ�5�`nl1?�鰭bkhI< ���0�����Ms#�>4�c�7�����8�{j���R@�o���$��;Y�|8'=B.'ӳT�n�hZ[�����	>�=GU�΁����u�@gt��mT]m�B��{a�j��(A����uś�ٲW�P���87�Q�(s2����>={ң iW^#;�2mT#��S���\�f����6�'ԟ��"rw ����ÅH��HdcQ�#7�hah�ߥ�t�_�I�Z��R�[��rx�ԩ�~��pI93�>?A#��,ׁPjg�Ѭѐ�YJ+C��F�nF�ќK�8�ڥ(n|YP5A�+�+.FH8y�n��%�6_HB���:�?�#��Q���&���x�����=2jv�V-G��\�8l����+�\`)�<.����x`MY�4s��i��On�V�	�j�i�C�N�̑\��+3	���7���CV���JP)K/�ׯQW
�H�KR>��Ug��ȜQ5Gc�z�s�tj�n�2��8�Ԉ��¶�T���J{����j{Q�X���vb�l0E1zY��tCL�onn�&І�[���I�1LN��M�������J��`���o�4Qݗ��(����^���Cr&�����������C�!P�3P�u��uX�Ӵ����I$��S8o��K�D�,�ڛ�-;le9�'�}_)�;�&huJ�x. i��O�����ťI��J��xw��0V�/Pପ��z.�z�ʺ��"<]�}�􏛜�/h ��c6��Nu�J�h��(xI8�I����MK����/��{w|�����ਞN�!���[y[,z��+.sd���T��%�N�yE�!q��}�ZNE����D�^�.�ٚ�55x8��	'���ɕ_'�nHp�*��cN�쫋�j.̡��7����	�У\u�����a���P�즔0v���{ō�y��o��[{������wù����ٸ/�۟��͓I4 �x����i��ߖ��Z(�μ
���c�'��=i���f[n�:0.�*�ѭ�~�O/�dM8����:�?�)��HI�'�[�P(���&�����d���Qk{�)�!X�,�@Y�GY\�J�Y,5@��GZ�����47���[C��ښ\���1H�Ge�Q��~�����`_�xx�3��*���g��Ŧ�Z�؏��%�dW7;LrH:��[�J���%gn�dD�N"��:��p��n�K�Eji$�\h(hf���ʍ�#��,��ޠ��s��$e�)uuq���]�<uԮ��,�3ԐFչ'�5=��8���RIP��hHmK���!�H�+2Y�xV�6��k�u�M̎�]����/�%%"'���������O?�$�o'��>"�-�;��Ƅ���ؚ����?l�*�lM]�7���2�{�����Ѐ�����rs@�|�ԕb['���,9MA��k��B��Rf9~i�*a[���g�}��M����2<�JALv����Jr�þ��FV���`��a�����@f3��'�l�Z�͖r��ȓ�"�ϩO9θJ�4�i�`ܐ�0�L��bṪfl-��F^P!Mk��w�F�Y�����m=~�B�����rAc�گ&� �oB�P����s�͈�5_hN�5��8qu\,b����p�1#v�X�{�\�KWm��t��r����R*(���^��f �X�|�S*V$��sex�cg���B@MA�^�B�F��e;k+�afb~���bC ������)�K�C��9�h��������.�QG5�r��<��y�zw��A�lZ7�t��C����=v_Z����P�{s\�E2 ��3o���ܹ���1񒁢��oQ�Ld�ՠ��}�ܴ,<E�V��� ��2��pj��yM���8��`���Q&�	's��.��[��c2�.�SstSk���t�3)`�8�(2;#B��F�ѣJ��`�YF��`M�J/ܒҲ�n���HP��	v��
��}e�A!�[Y��������i�Gȱ~@V���4C�;���^Qi!��fr��Z�筎
q9`R"��~��0-��#}��z��/�(Rdb~H��-��d-=I�`�^�yE1 B-0��H`p��_�o�3��$�.��w�ڠsWK#�����v���Tyt��9����ጕ��h�&$|p<xRIҦ��>�?Ț���hK�i�U��2ƵI�� ��|/-�Sϱ+�[!�dB/�᷑f�������v�e��*�L�TsY�q���ۊ� � �Z���2���(
A擒!���g�w$Q�����͊//�j��w�o��sTI��/Hq̨�3�iR|?�筺��iT������!��,I!�p5���Q�6f�U-@�j*��Q�(7�U��5�7������\�z�2����Ė�$�c�'��%`�&�TۛeP��%V��v��m�&_1L�R��_�[;��fڎ�����z��/��X�*�&�_g&�,����l4M��ݪ
,Lp�(6��,�B��ᄥ�o�I��s�L�K��ݴQ�ds�\@�<��n�~���l���,��|Ћ��u���	'ex�2�g4�/}~tkEa���̪T���)/"�� s�?{O�\�$V�*eC^��T���Ô������:�U6�\�G�Wd:�&�ϯŷv���/xZM���Z��!�����{ڦ��19({*�pH���!l�|�msZ��D���h �ǡܴ�8!j�$ғ���fS&i/���Ez���?��'�<1{�"菎��'
g�zӿ��3ԫ�5>Q�N��4y�gr5Ke�䀴�<C�u1 :/�h����S�z뭳������+7O�D�g+�/��$zW�Ĕ�_�TA���a>�Yڐ�Sf?q���!'#vX(a?>�'�۹��enSuQG��s3i�W�pPȮ�y�Jb�1$�������w@0��I���7D��u��!ql
k��]�4Z�Z2ݲ�^�����kmX ��I�m� �&_o4_2��o1x�B�Y+ư��i|/g�ʇ"�oC�{x(O�y^Y [j{�˻��4�r;��OB�^Uo�LdY}���茴?�&����o�lJ��_��A^ZB+i�v�XBA[������V����~�<���Z�h����n+����D��Ұ���sº[~�9Ld�%�HŻ�ԓ����o�{V�P�~0�f��j;6��oU&��)�8[e�UO%���ݐϜ��B��'C�Ƭ{�1}�l�����.�k�������3�b.QK�|�H���}�e�{���H�t�P��B��L�Ha��¹�e�JÂ�2y��kN�l���b�A�Å(�;�}�$�V�~)E���N�?܃R���א[Ix���L 9f^$��v�t�A��	 j;���Յ���
�G3����������'䲩�f�{��;�֚0�m�����./&�a4+*R!����+�����l�Pt��ȚQ㫤�Fg0�C�R��R�N$R[��t����ɗ��t4GL��x����dʾ툉Z�3E�=�|�����ڔ-8̑�-y~f)J!6R���<��ќ)���GG�5,����w�5�IW�#s' �$�m��;Mj��i���-�bR��b�B����kT�7����ّ��g;�<1�j��~��Yf��]d�so�C�*��Z�0ŀ�g?�͏��T��W�Z��?�Y`�RhA&�y�}�g.Z2�����s��*��_
����V�E�ط��3sq�>
u�Y���JT��N4o�������m`Z�}A-= Es!���oe��ZNO��t��iTY�5�AsJ�]w���m��S��wC,&���*L�C�$��%5��)>��֎vx�Z�b�U�1�>;��FK)���0\�N^��J��Y�1'�GY�pX�ح�13�/�i�k�+N�ϓB��'�����%޵��{��l�V��/L�6�O�&�+5�A��|�B����9-3d�h g*��%Ⓙ�o�r�#[��'� vyy`>4�1�6s%�}\C��a���<�����-�3h����'��]sh�Ğ���a_�IbZVrK|!�����z(��k��;[�������'�hP$p��/:���3�N�}�=�[�$��?��s�����R��!^��t�[>;V�c�K����I�R�"��t�]#���o���Wc�ߚ�J�籂��+�9�x�\��ceB��)"D���2��m}��V
I���๙��o�5��K���|s��;5d���I;�I4���ӱ��$+gU�c0�Jb����c�d�K��J�z��q)�z����Ze��!b�z�向�^��hɺt�O�[�w���5���n�c-��� ^���;L��>]��Rs^���3eً)?�k�c����ծ_O�Kf�acYN~vB�K'��UGUK��n%�@_��H�:���9F5���? ��OӯG��x��2s���I�ƃWҕ�g�O[�ͯ�zU����ڃHeȦT�LG1(P��cO���Ye*��&��.�V^k���
�N��K�����|��3�����ψi��?P~�������@�
�W$0��� � �U���sy�bЦQTV?�7临�C%�Ea͗�jZ�p�vO��#��
!���(Oj���M�����6n��a��%�J��omO�Js6����I！"�&: �7��]��HN:q̓��k��y:�#Xa��҇yPMK�>yl0�>tUR�W-��Ja�ykJ3�!g���%֥a11���?�u�����|8���j����+sq������NC�uE[��:�t�cx�{��P0>*�y�"(�ü�Ks֨^O����[a���
��h���_b�����@M�E同�bE��?ӒIDa�	��KZk�#��)(`a���aJ�;�;��Դ�V'�b��p������"�o��)��(�)�u�&I���tZyȩ���� E��T� �sb'��*�׷��#j6m�a���EP�������S9vK5��Yo�*�,xy$����A�����\�b�9�s�Nhp�fL����_��&p����O�1�[�t�hK�IE����9�K�vo�s��f�%S��������q'��l/Ö5�0��)I��$8����<�]1��"��ǔ̹1<�(�� ��!��������	*�gV"۱C8&[:�PZ^-��♊ڲ�F
\>�9�Y�Ԯ>4�#Uޞ���wG��i:?ϖ�έV�)�^�'{Ț�q�_c��}W�T7H>��!�(�^�MT&�o@|�+'��=�pU5�e�Y�gt��.�Q�cp�梗2�.5?{aO����ІfF�b����t��
l.H���|ObB �� ����C�פ�bݬ�������޶ݰqu�,eH��Y�R��J���Qjm$�s��Z,MB-[A�ٳ�W���o�]�1a�۳��6���\��K����������n|l��w������>�2.M ��������J��I@�_�l�L�ÃثUW��1�[ѽ���М��jHd!���h��О��rm׎cK��c�$I�nʈ2��ġ�=�����"��' `�zOn�BהѨS����8�=���h�Q�Jt��O�9y������gK��_�˄��LmϪ�_���I`'��� ����8�3���M� ��{-RE�Z�Q*k(�7�t�ī��m���rq���j�X=%��^���l�E�Ȏ�IoW�| ,���vz�Q��Ӯ�����@�u#�!�@��&�x�d��q�f�v`�XJ����x�9��=�裈0���o;���U[�)�R���*�g�U�����ã�
�η�Y���eܭ�ݬ�N+d�.t?�H.0��a�߻�{[���M���P�����/���M��Đ�v��������YΥͮ^��8{���bW�!!`<mG��h~�߯_��[�}���׏��ɩ������/�ҡ (h�d��-T�6_��Y��BrhؾDQ���WU�'�=������v��	������Aߓ�ܠ�*,Fj��l�5<9ZKc��<h���i�w��]Xv�N�����d�/;yb-i�w�*�|&[��jy������ m�� �	V�������5&�4P�5S��GE���J�wW���w�,f��4�j�՟E#�9�Qg�I�jY8U���F���=��$��h��a�n�ܝ[�l���H�H�λ�����9��3��Q`::�'9&P�b��E�.'���,��l�5���KD��W�z�~1��5{ئ�yy���FM��-��-�����?BT�DQrx1_�h�g`���ų�¨��%ޒ1�=(Q�n��n�#`M2�k�⌌��L�����g&�+��\�S���f�nxQ�a3���2�f0ǽ4V����O8���{\MBs�`��'xgiޖ? ~j��[��5K_�v�u}"ʶ�'{64�g�~;�m"�^8:�7+q�s��$��'����&�V��P��Y�n	w��>��N���J��rż�ňJ���e���=�d���R^DE��(�r-�,=�ĥ����޿ܠY��*�p��̾�*  ��S����tČ�X2&���=�tJ����������#��|b��*�V���G������g]YƏ������"���uK7������L*�fN=�]�Y�T��7)_�S�F�
�^����#rl '"(3(������s�W����b~��UW��-��T��A�) ���ˣ�#SC��1�[9h �'����bu)wm>v��Ctq�rDV,���q�C�#!�Y��a��{j��%B&��cK���3;�0=��h� ��@%�;���lCX.���7�r:NU�t���m]9/�\����juf��'�rz�rki�Cp>�eQ�ЂM�GY5�<�ɗux<$�.�78eK3kwSU���!�H�ˠ���B��,�0�U�U@\/���z�ɂ�C��Kⷍ}��z�j���b4���l�⊒~fƒ�0��KTc^��q���*�3��� #�`~�xF-Һ�����6���s�+��[�c�����<���mJ�&Yr�t�~]j�8�<n̢]�3�9��b29RȀ�a�ڍ ����$KxF�����~�;�E��=X,0~lH�;�5��
�\�8{6�e����C�_zp?�{C��w�G�F����t%һ�0:��vb�1�ܦ�B�2�º�Ft�hc�]]4%��gͨ�[�vn���geD�sa3z�5ƍZ�&�))�C�݌g�`��8j�}��qK��"^����3�꺍�6��|�m(n�?����B�}��E�����\���\0x]���P]a�-��y���5K%ttO�M��/��d�>+��"�)H]��S~�6@6t��X��SB�\V4USZ�Z���uGɠ&���k�5�C�M�`�����A��q=r?6JD�7��x�~2Nuxƌ�щ)����
�j+����dB�w,Ɖ&|66�i8;��N�
FMb��q�΋(���u�zo~�b�j�����0�\5�ؖW<��}��<�\���0�"�������ŶA6�Z{��/χ���{*	3�MYn.�l�z&�z"�Ǹ�S�P-�AW��4�y�@_|7n�8���s�إ4&���^�.�j�<6Hn���U�:7�K��$ՅvNFf��L)�Ȝ΢��Z�e��^zrк���_wZ�9���gL���~#��y�i���:ʝ'gY���˒��%#��בx�ìj�����nGx~wf?^����/�]�?��)��g%p�	=��K`u`z����C=�J����M�Q�j��#���[�W��ֱ�� �fUx_ރ��d�N-S�>xz��bz|?[��};�z��x 3:����A}�����(���i{	��iQ@(3y�y������fި$���������G�&��U$��?C�1���-aNˉN@f]�P�W@4��N�~�ra^K:;p�蛢i�[A�=.��CmtZ+�B{Z���u�P�}L�MN����U��3v��@��b��l9��i�DV�-��?�~
�נ�^'S��U�<�+�$S�Ь��,h��N%r}�%=&:9��l�E,;{Tڢ
)�O)�R���kg�����$�N'���4,s��M�t�FO5g[�:�d.K��8�ّk�1�vY_�ܯ�A~�)�O7�lKP>x���%�]�<`-:���N���D�5"�8��kay|E�]�=���A��?�г���Z�{5��,<�veY�ڀêE��f����xZ`�'�D�����j:n���dw���3�4�z�}:Q�l&u��cJ�|��{S*3M �*�;�/�.S����)�l!�'��	��]�{yn y��!ZL��$�U�X�$����d{��cO}	��'�&�:
����y[��_n�#�r�c��Zn%��o�}��x��T�����;�rnܑ���At,�/b�_ �Zh��:|��4�Hr��7w1y�(�'?��N�z"EV�C�����fB���I����i���E�p��"?"z�g��:��;�O��*07��ԑ>\������H���܊�[�7iD#��g$!QJW�Q��)敗��/N�oUq�:7�z��p����F�L�} FG�[y�Nh}Op�vM�M>P%���MRU��L󄁨�9"�o�"y�eߒ�4��}}�_.XY���5��a�N��L����u  H��v�c�(��B-ۙ�25iV�P�`>^�<�߶iFi�n��2�m�eB���_�h�Ț�3�8�(q[P+ӰP���g���|V�Cpy���Řʹ)�)`�E�QB֙�g���T��^�$	yD�f�!!���R=���&�J�C6 �c,�؜�]��� ���i�W��:�KXÝ����D��wf1�ns[���"Ja98q��bVx�sY�(�u�wg#����K��glwg��!?N=AB
��֤��끽�=߉�ԙpT���C��K�;��Ʊ_]!��r��	m�"M��
�.��+�2�RgoE�l�E�3�9���@���[�p�ר}�Ť���j�ˡ�5�+4g�&%.�GKb��p0PCS&��Z�VH�Ί�,��� �y��0'�_d�j3�#�5D+X�)hI����ĲD�0��Ì�$ŗ6����7��,�斧��Z�8@{�=��n���-7Eto�v�E�3��D�+4�V�66�L�(�>�C�G�KM����S�Z�5)�nN�I��Uů�5����'Z�{:{�����e9]���~I�`>�*��o���7��L�Y��ɓb�:1O�:��vW�_�0Ω~_&L�x�vS���H�8����O60V�pD}_�Uf��h�M��	�c_e�?s����~'#�f �䧗��Z�Zy�`��Ե�7"���ᡬ��8Yo���Te���^�#���EǗwq�E�Yp�5?f���k��> ɖX{w�ʩ@
.�����h����byA���X밽j��jk����d��Z1�ڒt;��Q|1��Μ
[�ob,Z\M��Bpc�]�٫P�z�*e�)�2+�g�ܷ5�5�I6���'�J2%!��|����|��ʐ�X� ٺi�D����@����}?GSt×<�:u��='��/xK �Q��zz���|��4��d5�ڍ�پ�^��#A���e �,�eԄ���ju���=x�	a
c���s��
�����`T���)���uF�I,�1I��Y�|P�t�����<��Am��ar�t&�4���i�Y�3�9���O}R*K�sP�S�U��G��l�*w�Su'm2�E[����4"�)qu�:��na@��U17G�k �E�v���"8��z0��7����A�HKO��`0���XK��K�=1R60&��?.DOM�i�^�y(\jzB�S/�U�n�	����Q\�2�҆���|I�u|���ѿ'2(�kY��Gc[2w��<����>}�x��
P|��3B���^�0<*0�c��䉝��^b\������)2��a�J��m�6�rj1U.O���g�b�%���f�F�������gϢ�� �DB5�_�&�=������O�X�Ӟ(��̃��=�Y�Z��<�N;9��mB$�LOjP�V/� `�l7o�$���A�+����M�����z��Ӷ�t��|/�����?�I�%�#t�=�l�SL��w����0V�sE%F+�Z�m��'�xĆrj���S?N��3����cQF 1�3sD��(Ka�W@�j�q�/߮޷�Cl!v�	^�Ms�
�w׉�H�7�ȇW�t�{�H*B u*��ytZ��cYq�9[.L,�R.<U ��Ŏ���]��:S��y���<����E�=t�!�O�f����9g����e�U�i�=_[��W�g�=m<#�=yS��I��`��!~L�8L�"vo����}j2�nH	\��T��$�SD�{ث�X�UE䀬j��KtZ~ �x�"H���@�����c��W̊��J��<��񪡾�m�F����u�F���145])�#�:�[m<}�zo����bYd:��IةlC�~t�U�R����;�r���D��━�@�̎t�P���=�+����]-�9δ�_��Ӂt����Jt�Q�;��}���X��0�����T����ڕ�X��B3�{:�$@h:���'<xh�d��exČ���3�oF��J�������x���v�N�4�N��)1f?�a)��$��-P��?[�/uo�m����*p�cf�F�<�z��ͽc�B���B2�}ZK��k
ug	%sq||F�o���B;>�L�l<ʡV����ݒ�5�C��K��qݚ��!�L��}$���q.k����� /�u�}s�H�~5(Dҭ�_p�(w�y�&H�K�:ܽh����漅w2Kw��S��p��{>Y��rjk56�$7�Z9P*D��.�)_�1!�J+��C�K1Kg�;>T�"����x%�/]�-fu�,��(\u���߹�A;x���F���p&e�;ë�ȳɿ����+�����j'�A���N_ʃ妀�$�S��hU{�Os��l��7qV]��?�,Ƶ�Sa��L뗮�����aZ{��Lg�!����Qua��rؼf���\�lj�cPeb�4Y���NoQE��3 s	��"VQ�fK�%.�pݲ�����c���$�=��~� �PJ�]1R���e�4}����bm�k�kHg٦M=`���>����1N��D$t�  �+=��ٲ*Wq��.����І��3+3����}kH)n]��~�7��;)���s~�|��N��a{ƱQ�ݓ��si��R 9�:@�b��M1��P� �{�[���F���;BQ�8�`�[����41�^xU0��s����GgcU�D�|��6�h���V���ٕ�����6's�Q�b�l�Z,v����T���-��}����AR(�~��H����1s�h�=�6E��/���m���Ӌ�\��06i��M�a�tX�0���E)���������tyT���L����@2N���;@%��r�A�3�XL�z֪Ҽ6vɱZ�\pg�(Y�G�7	�
/6�>fC�	w�t��#h�?.u^��nB�s�	���)�˵oY����%RGz�6MJ�U�4?�C������%����Թ�B@_ꅤ4��*N�����q�B&��#�ij~?4���)IU�~m�\�M���L�T�jJ��b�=WLWmRC,̷�E�6��d�C�*s���^Ss��k7ly$�Z-�^�Q\�d;��%@ZY6��F{������]���M͆���ˬ���0���������f�p�����6����]sl��Œq�hP����D��u���`�Jhi��$?�<z��`�����!���y7~��ļ#>Ĉr����!�˝5-y��z�� ��p�������F����\�z0�/�'�u��gW�*��g��8Z�h�u�.�[��J�~��]_�&ψ���2	��w6�&IϮ�W��F�//h�la�5�FH�9�,npS�
�}sH�.�,��r샙=a��Bg/� 
a��\{�r#��9��F��_W*���)i�̻�p�b���|�!�
�Վ�:�vy�Ԫ���>V1(���qmUb���k@Jϲ�ϐ"�xZ�{b3�Z6�,�p7�Br��W8�{oG;��lN���UN6NP��N�G�C�'+����:�q���V�|
j�i�(�H|j2����'?�|CH����
�U����^�A�ȷ�RƤE@苣$��fR�B|����${�.7�d�*W�Yԟ�vi���ư��F�<��� 7&G5h5w�'4����i�Ti7�!<É��ɍ��p�b�C�I��{��/z߂�G&<^���&�����,,7�&���*TCB�ߢ.�Կ�7?y�ռ�W������\OAzX�<���2�g�Wȱ!�����D���r ��Si�d��r�����յ�@,���s\���\�yJ���M���������p�h@��bh9�h���sS�t��i���Jt/W/�Q��W�>�' �T�t�V�\t����йSf�5���|������O7i7~�:�	ӈР镾�j�Z�.c{ɱm���q��m%-?3٫�gh�o�h����&�ܰ3%��v8��t���H�r˕��w�N⵾:B�5j�]��3�f������M���,�6G5;M���0�ۖY�i�wPSs�2E�k3��FK�}�}���j��P��>�Cg�N���x��C����{099a�p�B$6��y�\n����:j��f�&�d�@��y%׆��q�ȘR�b���{s>7���?ۍA�.heG�y����o�x򋷘�w����Z�&f�1P;C�9���{CNo5�hED���ߠ���v�Ҭb���Q����?�O��M��F$�?&~A-�fI*H�h����f�����s�;	�����0�n�'�9��)L�$�6���O�>阩��9P��8m��pXnNO������l<K�1,�+�?��WM8���N� �>�^��V�s�J��[��l$.�~���{IT���(�Q��t7������s�����ǻaO�*���9^l�es=9�R���Æ�N@"~e�'�I���M������'eo���������-�̘�Է��ɖ�3�|4�j����b��pH1�>W��lğ�o�5b,���I�����~n9�<0�,�z[����J�(�GK����&�".8�ai�b3�N�'F�I~�K��t��o�$��{���l�< ��Ny�:�E���Xչ>�"A~������c���c�����yf�k��w*�4��֊U2��-��~b�j/->���S����ʋT�W Q���ԧ/��z�4��P���>�v[kP�q��^��7 洕J��#�JAm����#u9����d�&��W�h���Dc�(��Z5U+}�\����Bn��AS���.cތ�TtZ೦X���{u�[��>��P�@o��yu�[��G`QRsD�'����8&b�[�I��}�w+W��¨L�����S������ǚW��Yo6׾���o�w���N1]� jkF\eT��8i������-6+�R����Ū��;��@[��i�mF���)�F�K�{�eaxɾ��T@+p��:���>�2�x�����$��z�n�cJsr	�֍�n4�a�b��O�D�l�&��
fe�����%
��૸E9!��z�(��&����Y�ő�q%!E��1�дYZJ��(�4S��r�/��>�.<�P!��G���>&h爴7I��0��^�P���;	�.�h�8��]<��}�������A�(DΟ�D$�)�m�J��� ʼs��׿������M�[7>�B0C��\p���Hmڶ3��d'�i2����K ���d1bo���g� ^��DO�o�"��k�o�m�s�:Z���~7Z�H�V$E!�3���׃J��"�J0�F�m���e�C��WD3��	h�l���y�C���1J�Ux�#�+0�`�x3��Hr�@Ϭ5�$�p\nG^�$�*��vY��Oѓ鮢w��@��uv�`�
ǄU�ba��� wiE��k]�l����Ce�E����v�|���Ե B����e�D�M-��BAF�O�裁&��'����4n�����'�<p���_Ѝ�x ����W:�����늗���[��-t�㌵e����V`z�.]�u����93�(糄�F��b��(��!䪜��c}�up�3r�R�]��U�t(CՁg%$�f?[�<����k~���I�"�Ԫ�?�`J�LT�M�o{Oռ�,��Jݮ�0@Z��<~��a�,��m�"z�B�f��%=�YK�k���8��+f��#e�O�Ij�e'�G3���R@L=�j#����-��l�L}U_Sf��csy5g�JL��s��DV��7��(��8>���p
�ؘ`J�$�:c�6�5\�-�����Ǌ�(�D��ͽ)������n�4�c�ʝXE͝-al��h��-%n�Gܸh��m�2�`�K�o�������ZLE��~(��!0m��J�m?�(�B5ٛ�d�K˱+��3�M; γ�cy�"=r7��fe�m ���D���Eh�B��0��n@x3��~��"�h}��s��t��H����4i��;�� r��<{�\��'?O�9�yq�r�o��f�W�������n���C�m�����#nfhRDZG�ӀM�J�I����rZ�\���F8�ECU��`��i�54��iuuX.��M5d�~��K�6�}&�,�Y2%�νp�z���zZ.ȥvd���F)W�M=��R� -
�`wc����w��1�CyQT�yo��d�r�-3O�ւ{NdE�Ϡ"p����{a®��
^�>�}��&��e4�����2;����5���f1�͠��y�K B�H���(������F2;�y\Ill�V:
�G@W��ͣ�����X��
��c�4��`B	�ɴ$6G�͑[n5"��!7j����q^g0y�8��2�1��;{Քy�V��ݤ���aE7R�#�K��d���xMC�Jو�2J�\�M�"͝��{�&�&���m�Ux�L����W*l%�A�ޢ��4n'�N/�6ͬjn�� |@@��z�m�W69�-����c��
�y^����^XU]K��w:�j>�∬�"�i�9���P�-�c���#P�6(e@,
R��`އ������z�u ,a�X��%�8f�Ѻ�3^L�2�����m��+ <�~�����UPIΐX�a���~�G�e1��zF����=�5[��q�(�t�}�ѪX����J��Z��WbN�{X�	H�X�ʀ�ʍk��n���d������1a͋3s��(J'z��Ǉ�����,��k�~Rq�I�)���7J7��"��8���v�O��ŧ>O�\?sJ�_��D�s<n߅ʳ"��F��3�ޤ!<�7�u��8o(<�X���%�!X�)���}��٫�Nt�ً��7�ҷ���^a� ��E�}�s�����un(�ޒ��uG�Q���
��e��H��� ,��j��ř��i�+�(�..��0����~�0���%�o�J^����<���a�o�Oeo��vp�/wF� P�P�i��ی�15�a����&�S=�ocC�]�E6��՜��Li:��X�n�T�f���A4��V���e���v�*�@���	���x}��S�A>��y�ga�W�����?�'��]Y��4���S�V7�^�-�?d�}-ڸ�b����!q�s w����8ܽb�4���j8�Y��a�"x�h���Fdk�E��E�_�v,7aR`6fO�+I8� �0����B����$��I]�8E;;�%�	��K(��.
ʂE���q&���ݷ(�n4�)��9�xM�.�_��YMz���SBP1�y8k��,e5XDJ�U݋y K#f���<����%��Q���>h�}:04c���J3׊�~$Y���8�oϘ�}�!O�C�P=�U�D�+؄R���;r��"	9Wua�\�U�*������}bPn<s�MR�o-G��⃌/D��@����[���I�bDK�*�,��(N��%M�NrJ��H��
����QD�PY��F�N�;a�E���f�#i�@~9�H�=�)[M4L�nLIz<��=���A�@Y��f^���h�m?RE�����__$26K�ҫ����� �un�K��^�Z"_vI�����R�H��P8�]��+���a�=;��CJ{��hͰa�+��ĵ�b�Q��ݲRf+�����BE�����,��WNЃ�Z�	�H��ψ�ɳl!Rw	(���Gq�oU����nm��K�\�yEG9/��4���"cC�4#�N�j�2VfvBw���s�@
�@����W<���<��^#]
���������J�1ұ�4�R���]^zPp�mEQ�#I׉Ki��Q����od�ķ	W�V�Y��+
��+f�-�=p�2$��X�b�Q�2�c��f-����<���?X�q���Ⱦ�A�Kòl=�u��e�0<ց"�Ir��^���D&_O��\�ɰ�K�=�-����M�IL�� �/x[|��S7%n4P�J[xc�V�F2�0��Q�L�R�'S������S�^�E}�9���)ڦ� �}��>��L�J?�ˋ�^ѐfd̚�lWZ�Zy����:1��^0�Z?����	��������V��3'��N���ГQ��+ҷv��YcO_���zvWX���p�"�2��p���od�F����b����҄M��(�'�׻lm(���PM�;(�㩶��6���
�y6����39#vlq4��/� >�ϒ��yl�Pr�붅����<שּׂM���}�Ӟ�qQ�<@�G�����[�4p����ǄV;2����r_��zM+m�J攼��#"�1]5��([�sގ�0�l�V��~���t�ܹ$p�y��K��0�g��Zi�Iଧ1G��F��!�����m��@a�1-�ڤ���(�[14t��<��~Ru�O4�r�Oa��T��r�6�G�������Q��H ��a4Eq���Z���ؓL,��H�FUq��1�o_���-)c���HKb���>ʊ~�`�!؈�D@�"'���)����I�0��3�|k.�w��OU4z����J�"V�8%�,����ݢr���T��S��KA1b�v��������$|���ѩJ^�����F���c���'�oA����¬'���r�I�*g���߆��.�	2��̣�m
ϻ���ΐMڥ���'D��<�T�~/΀<�P��		�F.FH������-훒��RI���������n*h�^:$v_��#-�h�lvkY<l���Z�e�"�S^�|r��M{���g�R�Psۋ��tW��1���}��^I�362M�0v��R���}:�=)���'����:"��F�$�O�)k��m,����a�{j�U�7dc�9�g�Jc~�dBA��[������v��4�<��>�p;��m5��)�d �F>�}9Nj�9��6ؒ��zPq*��_'��`�f�Y�S�`�u���ü"d�)��g�*�su�k�<�F�X�W��Sɩ�*���������6�ð@*�E�SU���$�>���4u�}FMĽX��@nJ�6��R��n;0�^s�D�TH�����W��<�y9bb%��}�u(�T�@�I�B���K���ˈy��5�p�CF/��]��6F$b67��ckM�?i�Uv�>�Q��ǤCfd7 ��ç�|2sn���~����LXhI�ȍS#��n%|�$_��I�R�!qmw�Nt�{�hټ�� �E��[�w20�Q -9�}�p�<��,�q�%Z�|{a�(޵��C��n���<Ԛ��V�ǥ�B[����;!V���8Ub$�;U&�ީ±�����������H@��N��v�rۉX^1&1�����u�X@����:��+ĭ�['��ԣj��hr]�+N��m�!<q�Hd�ɷ�O3i_��_y�i�_��b��h��WnI��>�K���h��w��T���<,�95�vW��&-�����ȉ	��Ҁg�	G��x�|��$J���ցL�r�s^0=2.�fX�1����Eo	�t�@�$ѽ�+Y���>,��=���$v�������=}	��SӍ �W���r�i4�"vEQ�6�"��X?w�Zc5�����]C���MVP�'�K�����2��o@��jV� d�,�KKfJ�F��pJ,-��I.k�m�Z�S0`N"vT�}0G�R��X�vI;��[KS��?��Q���y�C�N�-��7D?$��B�qc.A���}��.R�>�f˄�Dj-���� ��h�CO�}�����1�S֌��Fˆ��C$�i�z���է���S8��jq��R��7���7Bs�;o���YS��j�.��c�~�ɰ�˽Gݲ�q�~�:>K,89�f,��0Lͨ�fi������1��Y/K�>�V��T)h������'��T�TO�DD�j���}�Hr��L��� �~S��7�k��J�"���I̒�Ϝ]��/�Vk�95ɿe���SBD,$��Glۂ�[:��y��j����[��M[�o��Ȝ�u�r��$
�\�>-���;�eR�)�!�.��~E �G��Ę�4����ʃz�e%�߲���T��B����|ɲЁ`v= �,U�^��@�X�TRɃ�N����]cDc�/�f��H���a=��k!@k�U���ā����?��\� Cq+E���/�m�`�=��lϻ��,�7��N��J�3s]!���,����"�W��&>�-,G���UĢ�fB;+̌u.F7���E�)����Z�<X�����諪��Zh2�]�����Ma���P(��k����/D�FLҍ��n[�Lx��^�"0��^�=�\1uI�%$*B*d+M[�6.�cs;:3��)D?�Z��a�@��;�+Į�E�$-?~$�U��t��W6혵\ӿc~q,S�țLR���*2�t�Җ�-���0_az0���.��0獊c�կZmI|��r��LD�9��]��]��	��.�G[�5`X�3���W��*��oVJ��=4Yw1��hd2a�{*�'�M:�A�����;���@��2�q)�۸�7/c�Q.���"w]P1�oƕ8����~#H?���9@�I�;l��^@�(A�k�D�k]���Dw���.�SA��k��*�^wgB�a;P�. Wսs�_o
K��L���d�򚯝��	1�<�f=��<��)��U�#-��Y5�{u<k�έ� �:{U���2��e����]�õ_��!V� �+T�0���]~�@���^�./���{U�P��|�{�w��C;�"�,դ�2���K.�l���&\�<�G�G8s��=7)�
.�X���O�Sŝ'tF�^�O�����i"(N�5I8���v��X������x|B�9���J=X����O�u�fxk	��术�g�n�d	��X+���9��T!҂�n�azf��Jr��-V�{���Ӻ�]
�T�BP� �:�&9�=�o}O@0�s��U�/[���A��,+4�z7��w�VZ"w���V��}X�<�-�%�։��U�7�Z���@�@�}�h{"�~�\�=e���smŞ��R;�U��#� S�Ш�2�{�o����]Cq`�O�^���l�T��
�W9�UMtK�n�BX�IT#9TV�,��&"}36�E���B\�rV���q_��\@]��:��U�[5Df��6����tZ6�h(EsQr8ʚ*��B"4��
��},X�;�7��7� nXk�3}���o���(I8 W���p��~����bC� 9"� �VTxU,����3B)�.M�����j�]	�ZF����Sa 8>{+r��{L��몐
�*~T��_`a�H*soE\�vr��ꉚRLԴ�A!�Va?�JCw��۽���D�`d�-��$�5�'�N[�t�9D��x���gp��2�z����l閏�'hbM��ɱQ��L]�f$��{e|�ukf��"l�{t�;��M2L�'�#_s`��ۣՅ�2��Rh3�/-���u�q�bL�_��	yӞ��އj#�yJ�;0Ci�3q��`�(�C��]���M���� |�ip�NW�^��􌡭N��@��lzQkϑ,˯���>]�6������:�0�T �;�v��w��ԝ�&��������2�:�l�}��n��ʨ;��;���y�1�8���Iqjv��>ҽ;XX-�3u��b3�+�₢�o�{�R�l+<�a���V)�=Ô4|�jpJSUeo�'�b��W��7�ȫ��HU���b��`�;���P,=�%c$�$���{�v����A���w?=�d/�6Z��#��]���SR��'n�fI�����,�0>qH��p*D�\�i�j��+�9���'��-?X�9�QY� 	?R��G�:�y7=>�oy�Kk��vx/�"n�/��S�� m�n�]:[p�B�N"�ų�ݣ����>	�~�yҠ0hT�膩��P*JX~PD�e� �RW�R��Q�\�n�ï���)���'�46�5�H������[���F��_�cX���+5lK����'����8�`�d$�[�iY�������� ��Y}�<��A�ox`�R���A����
�쬅��w�h��Qf���%g�$�d�#���P(��W���sh)4�GSPZ 툴�%�٠J<G_�䔔�����v�	��1�ƪ�=Bj�M̡��Èm��ӿ�c�O�-��:��H
�e�����X�i�XR籛?��o��򀍱�!$�;J;FlG'���شxc֋�rw�Gr� �ٯ̉;��Ī�D	���#=.��j
!� ę�"��f��ɞ�p�:}�P�&�>�|��ɫ�Մ�A�Y��,F@����N�z��Q��ͭ�[��%��)gsO�i?���5���|�CaJDeK���l�+
)w�@�1h*���<�.M�	˂��fLvʪ�0*w-sjD�:�/���� q����\O~.%��#����M�"�"o4R�H��n��D�y�K	��Q���:s���x�J�Ŧ�����.�4��i��
j��#�[m�Ϡi�a�Cc9rTvw�$�ly��m)�23�msZ>��J�N��{l��\\����6��5y�|�z�{Ɍ��WrE������n��ӄ"�+�T=ݵ�#�D��E������ ��Z�����	s���w��jH��p��sd�{6H�Xl���]���A£WZ	�T�C���;o*[GB��fH&|<���03�������FX��;#Y�Nb�ŉ�:n��Y�7,�@F�&`��V��w�s-/������8h��Ƈ1�o�b�*b��t.)y�W��r!g[�����t eW�׈(��m~X�	��Z��I�� Q�+v"�Xp��鑇�Vw�$x|���4^'��iE�p��e� 5��&/�|��Dī�����}��ot�֞"����nq��q�J���-�;�7Hk����hQx���ay�A�WK�V�)�@�?�h��������lg|d{��u�7��C��_�}ʒ�2h���B^�V޷Iq-���y�Gg�������{KK�{��d^F LL�9y�p��"�N��d	�,Wv���3�]}�
 2DQc4t�0I�<�ծ� ��2�?!yԟq)��R�>P�>D�L�=��}��+>㉋[_�4I��p�\D��rҮ% O>{9��t*T�p�(�t�+��W(�'�=1lc��9��Qq́bڑ/kǯcaG�
�9�F�)~u�xQ&�Ʒs+�u�T�d�c��8y��8��&�:���@�n��� �����K��H ~:o
�ͫ�lK���G��"Kc�\_���2��*�&D�'��`\p�3��w���Dh~�h krm\�:JI1O�Cq�U��*�5�	��X��˯�U�N��	�����������瞣X�S%�JI�*"�-	�Oئ韗��^��f�mx�od^v�gW^�ӟ��zf~h����{(t?����!�F����7-oJ]$�!L �Q�ua/����* N�<���9u ���e�N������()xd)��9~�?��u'����#�����-��<��-�1�!Xd1�U�(3�PB�J1V �{���F��.w�#p0�*H�@���M����D���b#r5��9���1P0L���nϯ���At��ٵ͢Mx�����Z��1�;-5m���3�;�Sߌ���?t���o��=�����SW/>�J�@������_�Q��NM���O'r��lW[��;��t��!�L��q�\�$�����8/|���s��xU���u�-ٴ�,��=�@���2�h�v�~c�+��=	#j|�%m���`�����겈q��"'~qXk�Q�羚����:BSx�PP����U�4?�;K�@�&k�+��E�Ѓ��o�1�0�t� �n��?�[h�Kw"4�׿�9ϋ��\R��jE�@��T��SA��&�}R�s��I��������u�6�<1\�㝄5��o�Cef�|��Y��=�����?=�+�j�$l�PP��Ҹϡ�Q��!��W3mT�w��}y>|ńZIZ��~����K�&%:~C���mD�{�N;����f*nHܴmW��<�|�z�bO4��g���
Aґf�އڬY�{jYv��"�,��Q����ʁ�9�;5���.���8J�vY�_يI �0���ō��َMp�C�|�u��٠��$����䗟.�N��U�8���쒹=r��_&.��wv���?<@��w/��*#Q��ѝZ�@m���O�ZJ�:����pP�V\S:z���'}�T6���~�!7�f1j����?�a��״LH�����n '{HBY���O�8L:�ī<���d��W��p=�V����>�=Q�#p~d����z�X@�־Y<��{�m�@�����#]h�f�?Kó3'��ƶ	���������k�}R�H��A����"P[��~�lK�yiF��N�Y'�.�̱�ɕO������Ë�c�EȄ��bk^v+�[Sk�N���<l+��xYZ�t�:�=|�/�:ir��pV@���jt߃��;�8-B���b�l���(?��[y{�TQ����W�֑��$�3���	j�Ni>_��A@9��g3��q���V'q>��Z�k&N\.:۸�[�$O]��f8��5{6�p������ ��A$pT�L4�.A��6P�kV�}Nw�
�\G��/��L��*�l�
B��&���Ƙ�H���15+�SRɾ��0��io�Ku��C�����W�$ŵ	��w������y=�<,��\d鎃G�	,��;6n�[WFy�XX��g�)+aYg���L;!j��\qEr#���#;��_���lɩ�LJ��l�J2��i�	��������r����d��br��������.�SڀQ�<R�O��&o�}R`c>��0C�3��ޏZ$����ˍ]f�������}�{�̃V���7�2�Ͱ8#D䆩�S��q��z>�*�[��|e3>�|��k^�V�&h�g���_��n�K�+|�>��w�p����س&l�_V�X5��:���6�O��{��,e*�_�sf��O2l��?-�Q����P��Շw{©�y�tz��x�i>��~�����9�:K�ꍓ��5���h�o�X�ź���+���қ�Y̑�m�9��$�r�~�Ȯ9����8�U{�v����� �����/���
��'�X?b�2b�~11�O(3.�[$3�_����F�q�b��m��Jc@&,$E��b�*��F�@�Q�?M��V��N<�q�a-Y��mkGK�A<�D�'�����(�zՅ��9��s�l�2{j��"�{�Ù"`��B�!b�Z�6Gaq1P77mK�~����4H���'I�B�M(<�%rX��(���EY�w�=քa���h�0�,�6G{!I,�� ��� 1�8�5��D��K<�w�A9��!H�H���Tʹ��c{����$\����q�0h�m�[���mdc��m!���aQ����讆�Oh�)Uo�ڔB��[��08LCs��J̡�ϦY�OnJ-oû&OdD��A��[�M1��Xkt�����U��V՞�}�
HU��+��^�4��_�ts�����n�����>	,%#��4��j�p��Ȥ��Q%S���x�gg��'�����I?8�O�1�k�׍ȓ��eF��>��V�P*���G�O7Kc��5�����t+}�|V<)f��P\�L����L����������̎�WI�**�x��|�~�Q����4bt7������_}\hEצ��L)U��tv�+�$|'��@�����N�⳰|�&��5d��"{puݢ�ZlK*W,N7���-!г^�m�R�T�Y����Ռ��e=:6P�((5%'�n6�EJ���cYc죰�#��}z��M�,��g�F0����0�:��#ыh��0�`�����̃�Ϗz�e�g���&uU6�~F���jI��������r��j�Bto�p�8/�d(oGP�����zϢ��r�o;-HI�
x�!���XA�ZC�:�EAH��0 C�i8�~�,��x� ��x��i&ՠ"W0kM��5f_n,[6�RF����x�ǭ�4���č(��de(II}��{KE�-:�]\R)xZV.b�͂s<��Ő�g@ZEwʪ��@2�o��}yS��ी���$A�5��4�{��A���[�+��[c��
�H����'��s6�}K����S]���I5��(q�M{��a�vIx�������/@��[�}C���bٿ+R�����1!�O�}�B�B�q��,6�NF����3?���d����b�F�6~��#P���JOC��?8ǉ5yuf��1��j��3&��N�E��D[���$u��V9'F*;�ZǼuJ�Uh�X18+H���a�����ظ��V�j+c�W߭2���z#3���w&�Q4���	9F�N�1�D�1c��7B������q,QhK+`sr}C�[P�����4M��T�v)�s��"�O$iӕ�}�X��#��L��,��<��"^�A
���6YTp��b�1 �D���;��ـ̽�:��[�X�I����IF�8ѵ1S�� ��6u'�H3"Κ�Gd��oY��`�E�Bx��@�3ݿ��/��G8C���l�N�=cnC�;�?���c�'Q<�SKq�R�y�o���p���!*�r�!h��VG�Ԑ6�x�l}bA�rt /�p��Y����1�y'�]���%�G���1�a�@�)���?�����h�?���.S"ym��E|�XZ����q4w�/�vx<n�k�Z��A�mI����I�������}��Ym| �j��]`����?(m�5·<J�*�*��~��U/���@%O��>-y���]���9U7v�gL���
<Y��L�#v��ʾ����3ߠ��M��QWZ*�@1��_��*BT�[��r��p� ���~p'.i�<��Wi��m�o�C��-9�N<&,�v9SO1.�	%�~U�������	�� ���j;V�2~I�غ�@�-qÙt�y�y~�D����]�kf_����,����*'�8ܵ�uƍx�Nn ��U+1���)�
�Z�)�|y�Z��
�u���so ����)���b��������{������A���R����(`sfV�l��3�E�w��lw�c,�P�����'␭JY�
��R@�t��3��f��^l!HAr�N`��S[[^;6���GqvM��e57J����߃�ud��fӷ��+�n��:� ���%�r���)5�V�t�e~�}�W�1�΃��7� �6�Jػ�ؑ �4�[i(������2�]7I/��_�7����@��~�P����i���]�豶Jv �����Nn�����?N��P(E_x�z;����c��h*1IǗ�(��H�U��b��p��Q�ћ��[mm�dP��H)}g���YR�{I�?̮`t�y!�4,H䠜�A��5K\�2k&�;n�Z��vāULfk�ξ����A��n~'6���8;��e�V�Iݛ�r��&Yguu
�T(�9B�(Y�`?t6w�b���E��-��H�0���0r~���U��}6�ZF�L����(�
 j�. ǅ�򯊔� �ajFH]�	�=����_���M�Lt�t��s�e�e��xg$���Y�K��8*'��y�X�I���0^�P�����4�ԁ\i��?�} ������
P��T
Aԋ��ñ�I޳f����v��a�v ywHU.�\� ��!� V�ih��X]�l���A����G:9�c�e/��i�a��I�~�A�+�ʋB�ݫ��[6����A�PmRJ?C�,�'U!x�#�`D���zPr�y��5SE��wyH:��߳. ���
�t> 5E�/<����6:�(�.��+�mc�8h%s*�:h�6^C1w�Sʱ6�幄ݶ��!�):wT6���!��"Rt8�΀�j��>�Z5�� R)��3 ��Ik�밑��4�Ϲ[���V�y�6ucQ�椻Zk��t�]D�����G����r�����@C�J�+�0P�XA��w� ��L�/�%�C�=??��w�Z��:L�v��r#���$�L�1畷~n\w��uPʖ�̭����yy;��';�#(�f�_"!�y$DЈ���0yr���|��BOW��_aP��(�P/4�א��8�|L�⦂M."񳂶�D^��̝|6���K����硒0�ڹ�ݞl�I!���_�J���}��-�qy��L�b)r?F�#��C%`>��תM�5�z^Z7	d���Y\��2&�>B��k>�K��B�1��4�����c�z�x�3PE�N�k��,�)���k�V3�_�[AH9�)[F��~�Ҍ����{��y;�Û)�q>�*�ԁ�ϙ{��ҡɩFL�
�-�"���g_�� �6[�9�n��2Kk�~#YmW���n��h ޽��ȥ�����u�<���3RQdm��<v��Bl���
���s%����J��f~mȏ��^S&����~=�a������3(���� Ϣ7������a|W�bx렌ҸDh)�D���u~k�Z�<�ST�-�rO�_یr�i���$b���~!6�����.g����;�ǫ�
��^ސ~� �f��G=�<#t���
��i��8�F�=��8���C/9��9��ܴP��&�4z(r�D�;V�U�j��
���7��^;_��GfJ�� *�퍿´�cJ}���d�.����XRrh9����y����I3u�'�#Z��;����5.�r�pV�s tE%i=l����c�sw<��Dh��ӅWk~ pl`�qv#m��:�^�o��	q�dN�Vܽi�S���bU&�`������&6���A���gpw�[�V���dy!���P6�� �d�Z��_��L<7�a (�`���ͮ��A_�ڊ�[}XA�y6?S���.e�0��[ �T���O@�]����+���J��� ���`a��6��J�Ӱ��;J/
�i��Z3ǉ�9�>�63�P�c���TK��	}Q^ڴ~�UKZ�O��p���՝d��Su׿>�ƒ0e�j�ց���&��\w�$�.�}!����]D�w�BW�����w/P_";,�*Z+��W���c1��>g�4��+_N��zS��C�B�����ff5q��4�,T��璝��/�VG��k���.��>r��$������V(U�g'��u)ev����8ἃ]�7��τ��1mn]�9�x�n2_�段�i�p��J�9��k.�q�>��q��g`�up��[�|
ڂ�K�i��{9���������e�p�pb��wڻ����@n�baS	��̻�̉�p��.��ͼ���	2�k;~�V%eQ2�}�,O[D�{�;��K�mS�u]\�[��֫I���^{.��@@d�L��< ��}����76�'h�c�T/g(��V�OD-|��YPt�$-ci(�#��
�����t���V5Y�$@�����Q��Z�z4�`_��=�6�H�;���0.\��&�����"ɳ�>���c.&ɢi��|��&F��/�f�1p9ք�9xI�sL�a%�%��ʓ�^�w�^��K��K�����zn#�+��.}DI���"��8��JD�-�Ԋ�Nvw32R�-��)�(>��}����6Jg@�gd��n�𛢊�D����!u/3�u:#��,��+Z��`�Q��Rb�Al�2,����,��5���9��v�R�
�jzK�,	=	i��Go�d��?�l�&=d/R~��q���e.�7t�-�uT��_��������O5)Y~�F�>����kB7��˖�vu���*wA�Z�5-���w!���X�н����b��1� �L�W�<@Ԋu-U���@%�ϋFX��~@t��,�����L�.���C5k�����{hKX!�u7O��@9�:��~������
��4Wp[n�k�Y��`���h	z��	�Hi�G?۰����#+����}�&��mc[��ͤIl,X�7�x��@�{Zf_��	�R���򨉦��\S��!e�{�3��"�������NqCuc��ٻ�4��ȼKc���H���H���%#�������<S�Hz0v_Eʟs��9p��nD��������.[���֟V[�P��z� %�(�'d%�5ehm��M�,91�]Z�a��ձ�5n�D�a&aȟ�غ"OX�C�m���Z(?,w���i6�*��F��4���p�mq��"�BW.cԑ��އ�bDЫ�j/[M�7}!���*�06,��N�T"P	�۹��(��=���W �[@�P���X���I ��b*�rc�5��vJ�D��7����3��m��z���Y{�hw#'T��u(�O�{�n"��u.�t[�3��nd}ߘ����@=>�����ᵓ���J���{~T��e���庖Pa�3c��(�1N��ǌ��ҸJ���x]�-����Tf�(+,3�qsu��SFWޤ�<t�.N zMO}�:�����M��.X����z��~��o�Lb��A�.,����~	��8]��+u]�q�ڭI)��R���������=\�v�W3�;�;A�ϧ����#Ԡ�ȋ�AJ�N�lnI6WqDΜ�L٥7��3��z�5�$��/+��]�*=�G�8��tퟝC�1�5_�����6��A�cQ�K�p�r�V�BY�QE���o�{(� E���E�c�H�~���(qz��y'��4��;�J΂sӺ5��S .R���:TX�O-J�Y�
��)�hC�a���UūH�7���+��9!����̮n�_�[0�=`��\{{ W.��ڭ�*ć����\�sw�(��p�u/^����J�+7� ������c�E�� 
��-~͛/o�����:�y?�����Eg��4C-R����ǭ́~ch��m��Wx�?љ�Zv0�y,�&�}Cl�/�Tc�����͍ک��c����mlRd��� +�y��@0M�(�C��	���_NS�E����&���6�����K��`7`���(*9[�h�n^eKj�~��c;�{J��2$����S���vx����iW#A�/5��yMϐ!���m���pW�_�Ə9����~����>��Ri�qz����:S��N��[k
��ɺd� �f�o��n��}y~%�������o�c�7'�0�|H�;�n�3�-��~�@O�����l׳Guğr�y뉟�l�g�� V��N�Y�z��B�JX���<F��~�p�y��Z��@u���U������fۧD���m_L
�Co%S�'>�.�Xg�5�W�� 7�$���"����C�'���ܽ{t��NB�	4����<+�P|�(赍^;S�)Mf���0JB�����)= 1{Asޏǡ*�Bݿ�ikT� �ȭ`�M�`�N�����.��U;-7G�#��^[lj}j�����]��v2@������,����ɘ��#�Fv��Ы8���S����L�rc�)�Dg�r������i���P=�chF�1��'�*�GN,.��u<(�b�Y��b[�`�,���,�%<��>~%��:רcH�Xj��l�N8�����������?R����'�^�L�X� ��eQ���-�zd�*�o�5���0�w�T�  �zi3��z(1[S��ݱ3��n�{��o����ݘw��y�	$gm�@YC~�9]F�y��+nTl����һ�v����굪1�d��<Q�jK-�զ<����rvf��^�״�hF�#�E�))G�}Y�*�����Q'T�4�h?���}o��e����>)���5�����L���&
�B�)���>qG��N����� sa���Qn�'I��}~�ͬ�u�ش�%G�7�5�_݀
97N�	.b�}wKgKg���S룻	�4�sX�v�f1b���[��ނ���bH��%�x�Չ��p�����-��ܷP��^)ˬ@^H�<N��2LJ�Cۼ��ì*D������7Q�o1Ϫj?_"���ń�ͪ�2ƥ5�
��8֑�/`�F�U �/��+�˾�fP<ÿ�e�(�EF��g�0f�8/�-���"�T���?���HH��j�D48��(N8>q�Y�F�o\y�51ɘ�k(�A�/)�����w
x�~rBz�ԗȍ�J"�~�Q��*�i�]�����.ׇ0��b2�����IH֒���)��#�	!��LR q��XtJ<��Y�(�Ee�%��=�λf��o)�B]͇�y�k	�FFD%5����BO�3��w*�ܭ������mYTIq2���m�p�y!�/��Do���.���(IA¶�����j>}��`&�{�3�m3{XO�����~�Q��S��R��b�#��R�\J�ɇ[�8��`��]�����G�iP��]�Wʲ���[=6s��_� ��|�I8HS!,���-�όޫe�s�lI��U�h���-m�3o�����X;�9 ��91�oy��jR�R8���-���y��
��g$m��_�g�3�01
-��?cH���AM��K�/P!�����~��%�0���.�s=��ܵ<$�l�菭�3��+m���^H�s�t��@���P��	�7�E����3���ؿ`d�P� \�ϣ�Ԧ��a0&�S�:�}�B(p�~����M\���i��48e�M�U���� 0����:��>!*��nWO�C�v���" ]��b]�8�1Dgax����%�0�����3O�ø�s��3�V[�
�nle_Q]���┣���9�GW��iGХ?$�<Tf�a�§Xw���4��I,H�k��,�e�0F��<��Z���D{;�"_�C[���7?����;���~�);�<�M�+�O��אD���>��c�jk:K�*Ϋ�Ҝ��瘹�qz��Zɂ$'!�l\��._�_� q�d�xk�&{��5�85'�l�o��ض���\W��y\�^\h��Vh�M4E@:Yy�2������Q��A�mB�\^�Rә�6 @8´.e��Ho�m�	a$QZ����0Ǎ��v5)*lR .M��TyJj��z�P�܉�U�ψ�8W��N?�]�%=ؖ��r�/��Er
�α��@v�=�?����b�r�gF��?g�r�,��4�*[6%a�����b�y�cӽQ�}��е���wrU��Ϗ��X?d�/�ߥ�Ӝ�3ɩ�h��ɼۏ�,˅_P3i&������8Z�����܂��� 
�V)H�u��:W�ُ{q�p5���fK�gm��z��51i���~3$hD�0?^�]FʔPL��Y�a!�t@�d��藕Td�b�q%���;l��`�1�s�"L���6��G=Gg���۷9�h	�u��GRH,�H��VAX�_m� ���l��a`����a"8����Ɖ:Bo�C�)u0澣�s*t:M��%Y6��;�2���-�Ϝ!^��[p.!L#��(k����*
m0���g7#馶��x�4��Vѣ�^<L�o���8�{�ҙ��cg�c�~�K���y��a���p���ɣ�1�z|D�e�#3�R��m�٬/��&�s���Rv���o���23�"!R����R�r4Q��"��|^�&"���	T��2��,Z\`Fv7�\��X����S|��"�^�+���������9�����+S����������V������Y٣#-. h*��r<��m�<U
ي�����G��-/��B�ٳY�Y��g�8�_��g4٥"e
���k�Nc, �J����0��!�t��}� ��iYt�u��N�{�-����EhmF�0챴��6�۩O-��7Ez-f�<����/M�4^ϴ�g��f�����\�&O�GQ�;��XU��DQ�@^t�U~Ɉ��
��G�~"L����h�âR%{�f���f�`�e���C]ד�I�4"0�e|�>Oy��H
����\������|r����O���AE��f�
a7�F��`4D���ioc74��Z�U��Ҳ���8<�ele��0�{XF̲���'��V�Q�����ϙSԻ��������2�-��E�\P0��:�'�vN�?"�!�K"��SM��#Yw��5�y#�<�n��XkN�Q���p{G��p�eP��z'�:���h�B��,���ZYPFiO3��So�i��r��r{��ϵID�\n��L��%�Ǐ�u`��h���u���<�4�"y��^�A��Gr9�T}z�PNF�0�A�Y4,zB~��Q��fK(U�L��ӫ����=w�̫zd \�JP�yf�B�z�^�-\�	�h뵙]����f]q�b�d��m�f��*�0���ȓ��%,�ȱ, X[�d��cM��.�~����k�g�JV�6�q�i����h�"i��'��]���W���Ivh;��s���Ҁy�u�<O�YB�,@����6Ẁ�,�HG�����!ْ�P��C.G�2�u �N�
�:���fD�?�6����w�`������zT��K,�6W�u�*�}��wL�75=ݛ�.%I�~�e�P��x�I> ��%'�]���I�'��ft��L�V���R�oTt�ׇ�!U���h�W�"����y�S�Z:��9bn��aЀZ��qpl��\|�bG�X(2�,)ѹqA$����u:�Z�� ;�l~�����R ��C3Ɓ��Լ��e1���b<�~�3W3n�w�yA�>t�^Q�͇�����vF���;W?�Q"j����5���&_��ͼ�]u���tğ����aI�(S4�����]H���[��R�9�|�|��3l��d	�mlLo�*���pt��M�V�Q��@c4���m�&o4��t�z6`��w�=�܋T	�sܷ��A/���8��3�s6�<�%����_P@P~'�9�v7����b�/*��2�kQx:<0,U�% ��*Z�a��(�V�
&�<V{�*+������8���S��f��t%۷7�8:�dj"PG�`��+>����S}���.�5�E����Ұ�QGl�)t�YNUw�����w����-�2 !F:<����B���/+!q�����D��8�<�)h ���U�bA��֮�'*�<�1�
�-�Qz܋?߃���7���X%��	$����4��1���������+��{�@Hu�>�-)Sx�*�0�� ~--SaB�i���/�"���sX5�1�aVZ�\Y����lđ뻐�h� �4���r�PՎ;"A2*�`x� �r4�sAa5쇲n���[��͉����DXo,�bݱO����B���M��T4u�]-7]�/_w�
�;����n�G]8I�I��?vX͜�ț��R��Ҡ�1�	���_�h����<�OҐFvu)s�G���Jl�羊}˨Nm��]&����F3���=$�RI��?��骨��)�L��R,���A���[��d�4��1s
C�a�i�Ĳ�e�V|�&�g<�"t��L�(�޴��({�q(�mp'��������]2��ל�G�6h�qj�g�Ia���޵�w=,�|�_�OD����g��_���R��,q�#�zg��4�E���.c%��]��'���T6�� �8_�wBQ�τ��� ��7m�pl�n��͊�9�*������K��;�V}�M�[�^��B�_y�%m�/M�Y5;�������	ݖ�@s'�G�Fc4oh`j|�%�F@!O�i$+Un���9���P�^��ͱ;+U[������Ϣ�7���Fio)Y �N�ܹ��~�B�;�U�ue��۬\z=��*��a]s_Ź9s���J���x�@(�����~�D��(o�cGT�{���o?>o�����#VL�=R7��e��X
,o�A������1��k���1r�{o��aB#��|�ZQ�C4�
[��Zr�٬��$�F{��P���E�M�NCU�qz<�U�4�z��nsc�!�۰�E?H���Q�*�	���\�)e��v���X ��{��|R6�)�W)T�A���� Z��\�nIu�RVTx�P�[6n����������*�7/ۊ~���ig�׈���յ���㳯}�D�b��������5����j��^�pȟj���0x���cX�N0�e>����b9>��ۆʨ�3���{g+�� �����n�B��M��'S�w�!�����W�ZbC(��D�$;ҫ���'�sE}4�cP���q�����};;�o�������༐AƷ�	
�p0HL����q*�O�YL@F�7���j��q�#��l]�������f�=�f���ݘ��^�܂P��	�
��j�A/��L�$��~��jYkpj�-k���u.�\��Ӿ>����tW�_�����1�MQ��r�m}.��?�.�o�d��^�ғl�À�2��f��ZqYg��q�|�+�!�m��|�
��ێ����C�F{N�%�I��0V��=Dw~q�@$ؙ�wY��!dSPf�e������C�����y�dlh&�}��_�CY����+Oa�I��h@��ܝ=}����k�Q�ޠt��r��Qatvh�������GAH%Q���t���o4���E�jZX�*i���_�EƔ�Ǽ��y ����4�D�xn8_�:�Ū��!����ߨl��j"�?$���dUJ�Q�v���/�e������<��;�z�l\���8�-�n��Ugo��
$1� Q�.�T5f<,�X�m�bZ���C��J?�����&X�H��މ�P�G�:���'���QR7L��;���\3\D�l̈́�ܐ�X$:�`il{���Vr�
��-P���7��4��"f'�QYL"w"�\�:�'���DN
͂&C��.,t2�kӷX��`� Xh�������5�#k�KM�zF�s��� �c�k]���ϒ�lpMOE��9���;��>�z$E��E��oj�c�M�D�L�(;�f.�f�ݭ.N��Vb���*aӜ-&�iLf}m/��X
c��})j������X�YO]�������CۻN�K}
�;}hc����ب;�z�ԗ�6>��c2�}�7�9-�TkvZ�[�T�m]+뻢��z!�9Ən��(�G��z�~X��@�ѯY�����k07���c���Jk�@e7�r�P�D�� ){�&�l'���`M��	ǟ4{�)�������VS�a��EDͳ4/E��$<�Pcj �:�֜�t�Óv��A�G����h�7ܬ��IB�� ����~�ކ�o�埕��6�%w��{4*{� OA�b������kR<`�xA����c땢火��׍���H7J/aN� D�ȓ)�ζ��ޮv�׵�T��7��&1DW��ϒ_ei0�M-��B���¥'����w:=7C��P�br������������|tl����W*J�g�!zpi/U�]Z� s���AYVvt�&^j'gK04A����ByU�P�T��ͭ>�mf�Z��M�k�)���}p�I�k8{�Mp���[��|v�����v9�:g�[^½����_LTv��1V�
A��*��Iڿk��w� å�n3���s��b�~� }$ڋs�s�jT����'G��Q��a�z���I�: �3?*֥���kc-�� �6K�mHh����R�<���Q�,��4R$}1@��n�k^�f�L��j�R��?:wb�;"k:���+Ѷ5W<z�&S�1C��!��5����+�P0�з�| ���o��-�wG j#��0�9a��㿉ܚc4Y��e��a�}z�?߫^�pA�g�\A�&�����G���C)!K��%���5)��W��жؙ�O ��_Mrh�	�j� ��"�\Y�<�{�����P,��8��,=����D���]���^�^z�6�8��&Ӿ��}G����^���*��B��YĽD��ڐ>�Ƿ5���Ƅ?�l�I���F�F+�,�:6'u2���3m+�.��݈��^I�px�|+�����4�!:G��M�e�ն%;{ �g~�_��c�:(�X�kIZZT	��H� /�G�bϏ�x��`:m:4�,�h�ӮzM���xNW��G:�%�5m����&�����l-�B�����Q\K��"�.[����NB�ZU�8����f�Ѣo�a�$���?c��H�!R��u~m���c�$�h�eUʫ
y^N?Q�ϸ/��b�^U|��g��Y@���m��\�0�B�w�E��R���Ŷ��=���L�i�Ů���9C�SVI��>LŌs���>��'�_(�:����V��XCH���2�[0������#��Viy�cI1� �g�~)�En�m!YW+;S����s{N�&�95=o��ވJ�zU](M����}�J�T��2��x�i��ĸ�(��X�-�|o���K/n�f���=�R���i��Nx
�e�E���.f���^�ה���ՍO�"�^�k�2us�d���|�á}4Fjጤv�n�Rv��o����U����Ƒ�.�TH���2d�MYsƖ�:9�i�C���N�T�L�H��b�:b]�TH���		����,WN���'��[�Ql�4_�pq�F��/�,��"S�Vr��Y!�d�g��̵z,�.y�q�lE�-���~��m˱���螳5�`���>�0d�~r<h���U�5�
O�}�E��^%~nrO�=�\��6���("Y��kl�̉z�
+�7C\��93BR�Bə<p]�������ނ��2�y���������̥x>���x�RQ&�h�F��)��[����{F�g��}�B*������VJ]+\p���(�u�J[nD6$��,�MG�I�AK19~��:��_�C��0�O}r&�-�֔�F	�)ٻ*$���T���FH#��Ȭ��®u4!!��D|�AW��8ú�C�K��.���@�	��	���U��b��(�O���s^�ì����3�3fǦ�^,�,�U��PĹ��p9��e�53x<�@��Z!��NJ����wI�B_�	���������;2`���s��V�Y�n���<yG���D��c�r՚��$���Vz&;*���8��?�U'��ܜ�%9���P�U��rh~7�����ii�#��g\f��-�Q�Ól��p���/�?!q_��� �?��p��6��R#y%<�O���+VN�"ͽ�KKxu��d��oe��ف���W$�@�;��[�9w����2�l����HF"��{�#q��86�&S�G���%��"�����F@������g��~�7��y�0�L)�������,��&�~nor�I$��0��H���������1K�\ i������v��k
�-�/M�ɩ�3/��sǹ�h��0 �	Tea���z�m��.�n\�w
�����_���i��
s��ew�,�Z���'"�ŋ�(�*�����p�C��=��e2��5�D5�ݪ�33����C�ۿܗ����������<�0uUԏ��p��_�u��z+?7����L�ZhډLDZ=j�Ɍ�)(�j:��e�kfȵ���h��5}l�3h����rB#�`c#7x��"bI���SU�RBrc��NR��a��}ڽz�6�c[��]D�D���4�0���B�f���-�R�x�'G�� �`z�w�c�}V��+b��N��,�Bw]B�f��@��-P��O}�p$����S����𤽍�/�}����(�h��A�,;�Q�3b�b�⟛�-��C]��8���Aβ���-g�Y�0t�����ܧ�-��^*�v���z�h/��/P^c/ǚ������W |�����4Ǫ)� ���(��V�!��@��
�Q釰�u�--֬x&E����`Շ�q_�^G�6�p[�T.Z���g�x��N�$8.���M	D��lq5�9~���2��[f�0a���Ք�+:9�9�|Ժ9��֧�7W���'���WLw�����R?Y��;�����L>D��I�m�W?9���7��_i��:��p���lCP4ǀ��X]8�b@���Z�:�%.bu����ȫ�կ��^OQ�"6�����ØgXR�_>�����<�meo��|dL`��Ky�G�w�`�ˑx��K5����������H��>�S��NI�g�2�RZGo�}hϠ��8¹�I�>b�B<(�q	����C۞��j	�^���'��=9fu���G"Ж;�Y�p�<-����x"p1��>�T!�ZQ|/dړ�����ˆLb�$�-eQA��Ż�T����./=4k��v'��6��ˢ}�s�Dq�@6#;�ٱ���<�B�J��!�Xj��%$	j9q�I$�y��@�CK.��`����÷H]���i".D"wM2���"&ؘC�N)�g ��t� �?'@ҵ�~^���Y�Ŕ�G�5����Yv�X�Ȑ�y_���=���c��<.4�{�[����DD��܄g*T\k[�o҉p�MO^L��T�C�\.l��&DWf����\�e L6��,%�?� �D�IC!�R	����6�!�g��ۥTd���VA�7Y�n(,w���U� �ˬ��|���)߲�
��s�U��C���>�h�_�9)P��=$(4d���=���j�iw�"��G"��(�����M��E����@�|w~f����r��)�#���wDd;�t�hK�b�}g7ѩF�"���fRc`���z�rH9���v+�I|Wֈ�p�<nweY���f�8�q�UT��\[��Ru�g�ƾ�J����$Հ��
]:����Lxe<m[����fBȨs�&�O`K�x�}]��e<�`�Ml�_L��C���2��9"4H��;B�`-���j���U�V0X�+3���o79�[�sC�`O���d�z���g5 ������� ��E��4[d�B�>1^��A] &p]��,A�+k�|�t jcKA�,�'")��s�K��y%�T���qc�mPXʨ�Q��9l)#��ċV��BN/l����-������z��HΓï��s�,0}���]��s���u�+T������D�[�X]m��l��������w��|e'�Zd%�Q����Q᫾�H���Z �O�V��cS�⋜���,@�h����R,����g"C�Ȓ�)8���wl&��́�������X-3Q"�dC�\���ű�����0�i*�3^6Q����d��Gl�Ct`��#Z����Oq��s��rnț�'�mR� ��Yb'���B�CG�q�_���;Q�G��&ɑ3�bnQd�v�D�)�ӻn�������)�g�X�df���n,��~�@������_�wl�%��@���/�����Hq���fH����f;
�u��k�����(�I6�Cs���7��շ�E�����+����]�����{^T�k���7������!�zĈ�H"���h�h��y�༈p�ݽ�XUU�g+t�߀��Gu߻��}4��w�K���;=N��3�\J�����IM�~:�L�߆�T�HruS>��sXV��$�8?B>�ŵ�) +�0�@	3�z=y���Ӑ��8@�c�2���W܄v甀���t��u+�<�cTe����Zkl�ă����0c{/�PC2l����j;El������`y��ZYJ� �� ��eoN(x�͡�`�zJp�h�&U�JacޚW(�����)Z�|~&$�a`��c�E�����E�˒�m��|$o�	{�/�q�z[�&�M�z���\���%!�,GI�>�0G�7���s���e�M
�X=Ik�5���
rj�U��91@��m`]$���H��?�o�v,�z����cx�x�q[39[���e��ŌA]☡x�r.�חO,���'���\�0;6��!NW��5v�h�p��`^�ܮ;��'�Ia/�d	�.�-��8k�	"����A w-���IuMɆ��/���Pb�}����>8�`�gƎ�%�HW��|RX�UdH�.��K�		c��o����6|�G�?3v=4�ه&n'�
��H�Y&�@W��C�p.��hx��E��-o�lgQa��#�R��5,�Ĉ��Œ�4�$[���_�Z��>3+��!�� ����kEKw|QYS�{.�)�̶H�\gqTk�Bw��_Z�
��ٴy�jG������ʤ.l�-n\"2VA�(*��E�c�	{iP8�Ɲ�崵�Zl)��b���l¤*�T����i�]2����<@��?�5A�ھ�������t\��jq�Ϣ"���b��w=�h���DH�� w�n�#n�ΚS*�>eP��@>����ӌ%�)E{��Z�]��t�ho��%�U�ZU��g�*s}���FR�R��V���
O���ȫ�//:�Ѭ� E$R�~?*�B�h��W�a�F�~<pW�r� x6�{4�A��Is 柾R�]a��V�w�=�b~����y-gh���}�ӿ��榬n��Hـ����}���b�� P���Bg�m�%c*��s5�.)ͣ��r�#@��=�q�Sz
��Q�T�l��E1.c�\�q&[����Yj�91S0Z���'�&���y�c+�L�|���n�Nac����ҘO�$8��L��G�YT��ۅZߍ?���w�ߟ7�A�o_�k2<�q���|^?7�2���ۍ��+B|h%/H`X8�{�����=���Y��_�)�)1.� #¡����G58)t�L�I�n��qR�X̶͞���n����ᵝ���n�=��#E��_�	f'�ޯ�4ݠz�Q;g�Rח*X�1[�>�<�!tP����ةÚ;��&�kZ�~|KyM���O�=��j֭[�=^�=��ʈ���&�[���?e�7��J�F4�z%�X찿��`w�������óhi�����svw�q7�si���j@���C��;�}ϗ�^�!�S9��k������Q�lH�$��*,f����Hi0ǋ]9f�N}묇*��Čť����yf+��`D�4�d����#9*���cJD��u�a)D�L#�ܦB1|�h����D%��|}*�v��	1-�NVb8+0���[w�}v��
FÖ�>O�QU�J�rK !5�R�`�=��<�A�0Z�t��N�9&	��00\�4�_�l��J$��#�8/�=zM�Y���P�}�f&Uc��,n ^�T�߬�����5!r�CP�3��M�H��{���Gk�'U�
y�g�ru��5��Z����5�6u$g��"���lL��G���jC m�l�)�QvF����z>V���yWAU��<X�����r:g��=�x�)$��Y���5�����f��+,�PM�|3��5�����}���Q	���o g��16
��!k7`�5lYk*�F�1xd�-��?�h���U�RZ���	���n�$�´�J~ߖ��r�]�(�f����_���#�����z�T�$�֏ʄ�Vp2�������ѳ�u�v�DC���R����-,�<P֑��A�p'��t \�B�����Q�j�h;/묅V�`��_�%p��6�C��f��696��)��D$!�Fx�B}�7-��֛�`�.����M��-\�-GR�
4���^\�횉���]�C���S~
�g���{��~�S�1�b[a�$߶�_F]N��ik���" ��<�R����U�����T�ɯ6�E
��D[�����SQu��ʠ��O��(��Zt a��K��;˻�a�Q�·R��~c��cY0�/���0�$���p�rEG���Ñ�U��2*��E����Ӭ6P<?��
�$Zq�R��)�o���S�R	^�>o��,c��A��p*��J�!���f�*��{�ɫm��|�EK�W`��DI味�ԍ���c�qW�s��&D�e�h�]&F�+8���/a}nA�P�~���X2�>'���?��;XV����m�"�3�UA�o��/F�N��E
-)-m���A9�1��Y�cI�i���@2��mu��NL
�Z�*�;�c���*�(��/I�T}�pv\K�3��j��p���շ1���6�
��,���4z,WZE��Ь�wA[ҀEB�uµV��,^8�R�|�0���H��k�Q�&�s�R�$<�b����I�g�5��"��蔇g)��łٮ3ތ �_��}�ME��$���M뼍��!�k�{i:6E*~�����o�\/m'��zL}���@��2�8�[�
��u��&�d��'�w���΋2=e��&���Z��;�:v �\_B����������0��[Wm3��3�%�D*�O�Zhf��]��c2�43C��D6��`4'���u8[ۈ�_�܆��5�'^>�ڊ�*	z���1.�c�H�n���m�h�N��tWUL��p{�;J9trJk�}��t,��:3\(6\筝�~Y�XtX�:�YV�s6@j���=��bi+��ϾX�y(�*k�לgִh*�~/�Fp��Т��M�U��C���h7��Tl��9,ծq�I�d�혒��X>G��������KG�># ��5`&���:�x��Pĭ�Y�_+R�j`/�ͩ�pm�Kv��SU_���{�,�n�0����ě������=o���Y�=���:
�!�,x��2��I�[|�Si���:��u��%fE��g�� -�,e�dQy�Խ�x'tt;��!03q�	c�I��vK�9d{�Ŏ*4
'xI��-Pһ�	F[���=��ʈ>�%B"�;�7�n.+���*�ǺJ)���:4a�G���t?��6�X�8����go�V�	f��B�����l�oX�+�b�rĳPhX�{�%��G�!�tN��MlB}�Cs7d.���Z$�1t�\��Y��*�)����n�C�DI�e@)�j��1�G��݉0��7���
/�Fa?�?�j��\�LGo��_���'���k��-_�6iWq���a�2�~����*�x�-�`�8��Oa+@W`$�k���d��e8\��W��/�p���#+h.b^������(+�̖XX��5j�8@��0L��<�l>��If�\�e����;+ٚG���ӏ��S�\��z�$^����|�A�vN9Z��%yO�6ԄW俊������_<��;o�m�h>�@Ϻ֧	�R�nF����AQTC�)/��a�)�IF��F�iRJ�"WhI���t8�^�kY�r|�Y���58��|��������!ζһ���`�H	�.ם��+Q�LRm����j�f���"/X�� p�2y�nH���\D�!�y1lŭι��}f/�i3���v*c�f�7FL?���d6��6�#�(2�2�;`�\hCν�s���#��M� >�3vm�l�����p#�ok$\��bHw��u���r4!s�b�'䛫\��3����3�yx�ܥg��W�󠡔�ۯ�� ��D��!;�]�'��c�w�d�IwS.�3��7e����e�a�@��R��3�ZAx�D:#�p�wc��oW�JB���^ȥv�����ߊ��ltG�9[�\].b,�H���W܃@G�S�L�@��:�ڰ�p�O��sܷ��A)v���5�v���x��+�Q�p�,����G�-j�Y��S�����-�cV,"��!t��ͥ��[K��Eb���,MC$��O;4 ���"Q|#�fKǏգk�?,q65�+E ?%o(sS�����H=Bb��^��K	��z<:T�bYö��;��.�^�wϋJl+15wu�W�\r�\7ʫ�&;Q�6%�x,)��D�_U����(��E�H{���;��t��o
t[kOK+���x��w�m��-$'u,0�;\�{|�Saf��&�"ނL���B�ET-7�(v4���7��ֻr���y��b��G�����i��%�XZ�O�v�	��N��n�#_p�s���8���=�\��맒�����}L��P�f̋dNv����K��L�`��- +��$��mE�N�Kv�g�M5�5�\��~Ŭ�X�KG8�5L�F��L��F9�^��>�9��BZ��S�KZ�Q� �n�!��9�P����������V��#������K5�U��4��P�C�4%{�����7s�B��EӉq���G���B��Vb��;
�T�"y{���V2!����g��	�|�ϝ�ˉP���y�x�A���������Y�Z�뉏*=M�F�%Q�(;������"% =�~��������_I�k�ܾ�,�uE��bd>� �T��=�Ê| ��&?�(O�_�� Ϝ�H�_{_~��� �⼹0���@ƶ�4�Y��^�h'�]*Yyp�g�JP�7��e��	<^�&4h=k�%ׄ��7W�:SJ��:�(oW_��o��x��fO���u�snͬ�l����5��3�hྶ��F\��?h:�w�׉K��?n�
*�se����s ܊Z)6��c `~�y�-8FeM�BR����XSť��&��5}�b׶��V);��ѰHޛb�ł��@Ҩax�З���P�SKƥ�|<�{"QS��Bug[����fh"��2A�cU�k�񬙦˾�!�|�VO��-�v����)Y�����R�mDJ�������z�因eb� ��s��ߡpʽs��k�L��!���hp�}v7H��^*��}�S�)	�����r
�}���R�
��ւ7�*�z�h�*�xY��
��;�,q��J\���it���9N0a���;J�3}0\�TG��Dt{�YJ�8�{!���%�����O:.;�s�V��a~�X��+F��u�3��i ��|��ˉ���l[в���T�c�p"b�e��IQ0v5�������S�N��ǣ���w�>g9� �v��6y�g�Y#aG�� �l�l_Ub����~�7a��$#d��A$�]��v���/~��^�"��R����N�D$���6{	%��Y(1+M�Meb�C��a��Z1�̯N�����C㷮�ƥ�d�;>�\T����4���yH 9�x|FN���Qp�)8�h>M��Ln_�p1������p�_c%ר6�bcݩ�=`�ĶK(����b���[�4hi�=�#�>�ˌ5z�1�pN؟��%f�o��1U�:KWldv����#�#��*Z��|	��pw>��L�pK��ńTY��a�78���v/��NVV��P݌��eB���p#�GgT����;��6=����*�:��Q84p�|�B �6���s%�^���`E~��Nʫ��z��F�5i�o�򱜡�r|y�@���\�Ep�F��')�F�H�t;�p9Ѧ>�U-�*)� s�*S}~SO�m�Y5�_�(���Ϲrų!���.�f��q�$�J;�(?�5%� ��z�E;h��	L[������܇'�4�FL��Q7����a��[Xzh��18��>o��
�ª���?�0n�����)�*�M��|�T߯j5���;7���,�^�gy�qH���Ē���83��P[t@�hZ�a��u���G]�iw7���r�͵W�̫��aJPZ�ל�Qr�pO�Z)��"��?�X����F���vѹ{�5��g����/�Q������kw�ٷJ�����hq�yQE�߻d_�I�G��5�MYL�����eF��;�-a�_Z͂&g���w�<�#��7�Sto�ԋ�,��㡵IkbH/��Dob���e6g>j}�B�]�غ� �4���33ZUq��-ש�]�9&|*_�D�����o
�w���~O	���>�1�wAe�vWu���`MB%���c�3+
w�4��[��BRQ���d��T�˴f{]
���sɆ{��t��-�)������=_矻��S�V��Uf�@�_}@�j���������S�\���Fئ?�,����Ԇ����M�2|vU_&8އG���|�R��Ɍ\EM���g��Qձ�=���Vb�n��w�_�RL�/v�,��0�rߴ~�x6��(�.&�_ƌ�
��:�c�#���N�Bc!������*̢�F6������5M&��0'q�r�kݙ*��Q� ��W�>'�� T��ƞ˔[+K������kq���}U�tYS^Ä�tdBo���`vJ�ʳf0~B�0�D!(?�2P��4���<���hw��[�8�9غR�[W�cȹt�4��7IPu�A�O��� O{�{Q�VY���v�o��!�¶K8Z{)��2���K���̡Tc"bL�db��6�%���K�[�v��"`���e��W=�S�K�`�@�K���́��_�p�����
�=�M�$#я�-�n��{�Vh�'���o)��6�LVb�B%N(Ug �ƕy���E�_ݥ�>�b��� k��_���q��T2�2�"��G~G� ��w��� ��Xѵ����>"�#�N!��s[���յV�ޞ��OXW���9����ş\̨A$G^{⪀k�X�x�*��,)�v�F�@f쫲ŏ�aB�:�DО���1��-��m{M���5�Zo��B���G
�Z4!ӟ�E���l;���0��8
?�fJȬ$P�%�qt�D�\�?"e�Mَ��ca�X��v���-�Ô|�j�">�}x$���h/�ה)`��|�I+��1��Pl3D?�mZ�&�E�q_+_�Tl�~|������r��)O(K`^B�/���ϒoN������f`R(r�2�O�*��_B�ڈ�<�n˽���5�~: əG� e%�d�@j�TV�,bir��v�K�����Y*�X�^�z�X��Ͷ�F�{B��ߐvN��fA�׈��,�Q�TR�+����<�G�"�p��d1�:&8�0�2 2z���x����u�r���}��GO4t�%��k�S(O�Ψ�jt���Z��[������l���Vة�����,��N�i��P�%Ȗ��E`$/nY�y����lL��,D4��K���	J�]�2P�UE�'�4�Rt���o�}��:�չ�~>6!��Xp�T6� �dI{NcA���D�3�4s�!�=3���wl�>EgMk��� 3�����:E+��R�Q�/g�:�:���z�ި��}�@����xD�kz��K<kdn���t�������
O��k�^)v*Vֿ��q7V:��B%��Ȍ?�]8!��k���p�� R|����F��RK��^߅+:��h�����j������Cn�[�t���p��l�l��ϔP��f�"�r�-i�J����
���qr�?yk}217��}Om��!�ǒ�0��hdU�P�p5]�v��� d���(R02&�:��˜D�BBʲ�[*=����24����+�z��4�2u���K֟zAB	S8��;�"��f*�C����=��>vL�3%�WvZ�(
�q��!��c�G��8��X�MINN��eA����A�Wȃs̀B�ܣ|��h�־R��=_VB�(j^`2Z�^=�]���ڝ�G��}B��>�[%l�4�y��&����Oޛmf��(��gF�K�Z��w7�a�l�%�P7j2nK��l�
E6�Rs�F�]G��ΔF�L;КҸ{/͂J���U��F*g-iVl��i/����"��+�/w��k�;Q�W�$5
<6͹u�!��������e�o���e<l����37č%[s���瓓�ja�}(\R��O:��r��k�|�O相œ����=��D�?�>,��L�N�<վ~���Yb�F�5f[��h%+� 2�.�\4"*k!ڀ�kk¾���O��V�1��9 q��8w�m� "�� 7�}t��(/}*��`=�N��v���BfQg~�^P���G2��Myn�!����kC����O�E{~n�9f�K�W��k�]�9v�V���ؓ�%��$i�aGl
.�2��(��&�#��*���ඈ\.�]n�U�%�W�q�r^;3!�0�E�՝jʬe?��4�"���/�RLPs���{�2�9�k�Do�nAB�o68�ju z�I-���Y&\1+b�؆�����#�G��慏�vU�/��m��޿�}B��U5 ��9��m�����[��D��\0r����~-g�	���^��<�>�
\�3F�7����E��z40��*��o����]��i���sL�hL�C�+	�>��[�ܙ}rL��Ud��X:���6��N�������o�FF����) �9�$�F�RA5��x?�৒�m�O��D��J����v{Sø}aYs�u+M.~���z�Z��Dh�5ȗ��B�'�ʀ%iK|KP��&��2:�aFq��b�����L�^JBI	����Ca����s!
��e�:�RSn�	!�ٔeOܾWt��w�n˛��o�V\�h��G�}Wb^�y���*z� _e)����LVht�_h�� r�:|@5{��c/�P����w���[*oq�xG���pyeD��V��Y��韏���H�@�j�����0\G	S���z���������%�S���Q�-�Ȉ�v^��r1�n^�o7F ��~�5O, G,w�3�7�������&-L��djv����p4��P��
�[������sb*�
���L�9��)Ȉ(��ZH���n-}3��֋x��5�%ܝOƮM[������l��Pp2����6�e`K����F#�K|���,G�LG6�yw����bZ�>jE�?jn*�p��@m p�J>���Ġ��n@�r�Φ�P44���m�=��$��3ж�cRI�Mj��)��;�E�.�w�E���{��hk�OM��H4�'�Uk���Ň���ا��g	�ۣ����� �� \��9���;�:7�/Iԉ�����܂s�I����U��kp�u���1&j���>�o��%����r����_���vn�&X���6s�!���K�<��8fZ�3/0��%<���H���,��\1��~jh���V��@�_]���\����mb�H��w� �,s.�+����E��o���c�xnÜ��Մi'��1@���{�_����x�� ��}�u��Q&��b�m��?R�������d\����ޑ�9%�
��9T_�8���O��i(��YVv�F�EhF=c�-�����0fS@�F,������!=q4��������.�������iYͫ�}C��d?�2��p� ����B���gB�`�39V��ݎ�:�|����>w[�I�e�5�4Y��h�Lmf�\�܃ɹ{4�Ωr�Q��َ�"5�+t:L���YIǣ�E��<�T/��'R�����R�{*U�����褎��,���G�ċ����	�ߐ�O��O���� ^S�(������G�"�����>"�o�+2�=�Hte������������38̹�o���Õt���'Ԥ�_��b�	f���0��b��f�E��O�KM8�iҫ�SD�AvRV����ˈ(��^�X( ��aZb�$&K��(^-{����v�	֝w�շo똣�ι�xlmoUB�,OZK�3�^6
����Q:#λ'"=�F.`��x��dT�	���5�gu��I�<����@e����#9�l�e*k�(�L,O6��r:|�y��v�ya��1���%�m٤��<����=���'�6����~�T�\��f"#�KP�9�8D���uO찦��'x��24!a�QsK)��*R��_�1|A�I��}g����M������H���]T(T,��1<.�g��1҂�D��0#fFo9��q�Q����u�Kl�5��K�)���R�/��s���,��F�����=�,����J1�uq����G��(��dt�6�c
�I(21�P��KP?ޮ��)�dn��{N_�3��N��m0ja@��� �5��%�\������<� ����(�L�Z����/��+��D?{��0���e5uPn;��D�d���C�����0DsA�S⤎���e������̒�����Yd�e~׹�k��&��v=�l�)a-�15�+�Y���+O)����3�!AA��Jѧ7$?i�c�0�Om���/�P��<�g��N�$w�b�=Ea��<�s�/=�b��(h�H|�k���m�R,����o�*{�sˍP���сwƯD�U��1���<��ܗjϬ�S9��Dc�<w԰S^��n!�)���&L��/���r`��.cr�������r5�|�Y0U�8��%%ڃú-QOb�d��������S���+瓲���6�K;�H;�!��Z��H�/�M�2!�j\��p�ot��&�\��*
�4,nM0o��@&ܭ%<�H��Y;w����	�NөȉO-C��*��[��Z���������XDZ�N��%	G��L���y�(!����'� <_R���L��9�Ƣ�V�<.(N��l�KC0�z^�$�i㈩�ّ <�K�H���?`���#A�(�d�L�"	kf����kB���b��n�sA��'���������s�e�r�LkyE�2`zk�6�zɼ�N�I�<ͮ��&�c�TWq���*N���&֓z�����k�\�L���4槳�M���%�K�u>���ĉ�E�4<���i�[L�=�&V��E;�r�_��i�9��د!C\�����u<�1Ŗ��M˚�f6�※d�HM�,�58�ݱ��2p�G��]��l����:B�!VSB���ϻ�u�TL�e�V�C��[_����@ި��� H�^��V&�Jw�{�ǜ�O��?e�]ء���[ ����S�iUl��4�����������{�[�*����MhA�a�D�4�cܗ5rg(rC�øl����E�c�eoO-;���U���6����`{�K�}<��ѵ��r�0����qH�q������ʔ�c�]A�1�\���� ��bhG	6��U0�����l�;w�~ю�!��<A3�q�@��1~�I��;�M���0���;�~7qd0+:p�"A�u�J���q��gK}҈5o
(<+��TN��$��W34�#q��e,��v�7�-�".z@�xm�	�M�����0C6���k��?���Z?p{�N��-�Z7%��5_��2�7`��'��C�[������ъ����c_�� (�3�|��� z WD�z�i�5�.Ϣ@®`{��dQ+�@!�|��3I��N
�/id���e��j���`��z��A]�]��ҝ&=�s��!��S�i#�l_бO����9������ 9�}��M�{j�����r������*�c�gf메}���|/��|~���&j����P	��5�n�*.��o��s3wMf� I�ۨ|[��|�hUalm�D�玀����T�yӭ�r��@8�|�B���v�\��������/K��ieù��G�y�[X���@��$�;c]�^|V�E�}N%��i/�����?�s!������z0�D�P��SI��"�N� ��:u���	R�;�_Yw���s������~P1���T��+]�}z�f�J�HㄠDpZ�(�%84�o^�g�>��p��+�6޿�^�=���!�K�=;=3�L"ʗ�T"T�G�Bԡ�Q.&n�F�g��&�x�	(E�х<�(�Y��{%�x�u��
'fm��<�էs��Fr�ruܩ���|�هХ`�i������ʢ�-3�s��V�ZL�:�"=�$|^��m�͡����ԤrPR�^i�u�xR�h�|fs�2JN�k���v��w�CC�K p�~?���-tkYM=�H|@�M]&��r����{RLDv�G��5ɛ���X<��n?$q`��Bf\�_� Hu2g)�[��6~�w�*6�<?��4���K~���H(Ii�Na��F��\F����sv��n|��\ˮ��I=x�P�j&f8�$�m5�݁AϿ�9���WǦ���Ţ:r:�r��:��< �g�Q�������cȔ�a�갮� \�
]h�Rj�Q���7���<�V�((��P�а:S��)#$��}W��/^+��U��Q���qb+�;[����ݎ%6��([�}����R�;a��/Kns��r�i2K���@�>Ѵ�A$���B~k@�6�"̾m��;;2�T��7q��O���H��O�Z��%�D���(%�l��Y����tm�2�=�f0Q�t"$i���ޯ:hޞ��̪C����]���A`#%*�[�;e�k��������@o���	Ί�x���o�}j�Y)�݆s������dO�͘��G/���ata9��Fi�ڲ	�&�N�*1�&�Hk�\UK}�I:\�E�ШI��.Qi|��-���g0h�]�C3Rd�.�_�c!��d�5�ls5�i���
���������Qm�
��WX*�.��� �hOr=�1�<Y�\��u��X�}{��;[ht�\H���U�W��?�W�L��'�;�R����B�ģᴺ<`�t��k�wkR0�/q���'ݐ�v�R䉴ӧ�gOG��F�����m��ZJl/�tK/�\Q0����ܤ��f��Q`<z~��?�J�JF���jr�o}��'�z�&B18�^M���F���_yn
�We��y�O8=V�_��V��<��f�Mļ���!nX��MQ��Ɍ��T�:Q��,��:w���BD����UX�t�F��O�,M9`�Q9-?'��C�����_�5o�ikѿ4�3)�vl@�
`�(AQTb8��9��=6��((⽁�2��.늉�Q�0���-�s�G�"�(�4>ö��p��n�s�ο�D��f��jV�ޛ�u��fX�9�["eZ�jj�f��H�w9�$h�����-�*B�!-]#�`��mY�O�^1LvR$��t�7�d���׉���;l�DC��7)�Փ���������N�r;oq�ia5�b�Ig�ڱ���2J��nD�o8:ce��J�ce��Z�ŁS\݈.|���K8Nwt� �G���4���q�8[/i��EQ,c2�����<�cI��Zt9����[�o���ՉƝ-P�
��oQ� �k#����"=��+x$7ª��-����EnZ+�(�q!]�'�G����4Kz��T���5��>�ܶB�k|G��oX �(��F��M:��E���/�ֲI���-ޥ0�f�|���O����|6�g¹_�LF0����|�*F�M�K떸6�+Ķ{Z��������2�fK��Z}��j}�����Ӂ'в��s�h������/��K�m �8/�]bR����B�.k^2��9�y���+�cs%@�b|D�x[!VW��$��8���@�	N�`��H�~bo^����D�/P�� �>5�
��ws�<�p�ŉ�et/u��AsRDբ��(.<�2r�Q<��د۵$��-�+������k;h��C�������O�,�+�������k���,�EK��r
��ũ��.�b+o?�<�n��6{��+rkB/�r��y!yoY磰���(���5!�aB�Ҁ����%�X؅���.,$h��'�+1����b�)�c2�	FQ�
��gQ&b$��{�
�O/Y�ݭ�X�?�y6Eô�"��e_��>���#h'�Y�s>�~�ok���O>����bP�gs�F�D���6���~S�9M)�,�'�c�Ix+���ew�O���I(N��;�%0�G�{��~x������f>�(q4kmp�|�cN��2[և��\|v�'V�WM�gZ����!e_PT$�/��͋�D�'���5W|����ܐ)n����Kj�	����yw�1����>��0{����
 ����mA�#P�o9v,Xǐ���%�]e�%���'��U���\���.�_{~<a�,����p\�˪�G�U�[��Lf �E�_h.\�Kwe�&����ZC>�=\/�K|zu��<�A�5�l����=V<��E�i�X��m"�Z�d�(Agq�����������۾b�I�jWxr��bӌ���.�d'��Q�S{��Glf�F��G	�"%L,u�(j�!&�o�*ޜ ��U+�b����-����������@�}���g��Y�8_W6�ۖ�D�����κxu$W�<��<��J�Z]�d@M�^��f�jg�թ~��7߮�L6�wan��^D})w�ap):f=E�k�ǃO����Z�;Q�]הDJ������4l�<�c�d 7��T�PA�FL��FC��Kc�}�z�i��kڨ�����nl9��1f�&�\\��f$7�)��ED��e)z	�0I��3=*M�H'!�v̑���&g�&���
���~�)�Vu.�
�W-�X��yvI�&�1��r�<�Y�8{�?�b� -������|�嵗�����.k���Tz�r���ۺDzT�������f�_���*M��.����.Ow}���l���B��E�g�f1�N���E�Ó����`&�1��p��;rcD�_Df |��ꥦom��h�OO����N�W�k*��  nP��
��O�Hޯɷ����U�FX�V9	U�{�V'��8	P7�xC
�QX|�]U�=�,���ĺ�zd��Ro�i̗����`U� ܆81� (�Vq	�TM�`��}���}j�y�W� Η`=�(���>����� O�|�Prtt���W�6PT���L�Ϗ��R�m��{�|�
vJ5&W�>�QG~�����o��iLǡJ#pb|OYA��xә���?W�kh�zE�za{�{ֿf���UO��vv����@����h�[��>��g � ��F��B�'�ݴ,��ST��*��1h���=~��H���Սm�� �V�-��'��j�)S �^�n�����cgS���d�	�^Y�f�O�6��Z��^T����qQ[!� ����
����O���;v]����f���.�u��AL`G���QIΛB�K�`��:�X����C�1����k�YF*���Nq{�zWzu(D�cٴ���b��f3W���&2����#��P�D�Oю"p\D�B�"�~ҴcL��H�ᐙs�S=1��*v픉��Qe�E�P���v��*�*�*�<B��4�8�xiq|�5{p���G�K��`@J�1�K�v�B��9�XUolu�7�3�/6�.�LJX���=���\L0������*�~g\.����q��j���=׈��O��\[h�5��w$��u��.P `f�P@�x���X,H� ��}ԆbQ�y�Z�O�UG���LD@Nn�X�Kd������ڹS�܇��N �6��^�������A�H4d^�D�f�߄���0�qt�s�]�IV������K��UP�RÌ�c�Po%��h�!ұ�g�� �yc@D����/'$OX!uX)�,eN}����e,i�]��l|�{�FI�����h/���)St�L�x��|I�Y�w�(�bx5<�\@к���{�#��9���%J^��^�[RF�� vC��J�ۖ6�vܚ����_�7��9}��k�Q�J�M��Z6=+�w�v	�\�o�!�6%%�}��MGgJ+lЀŷ�����Q�H&<��������e=5'�(X�솅v2�*<@�EW���V�C�_�N"KMQb�� ]`�|��s� �c�c�,H'Q>,�A0�?}��w��P��h�wx��!X.�I����] �{��L��<_��i�b���\��<]����4�#oj.�%.�^��U�(B����j�����(���`0.��_�)]O]u�<P�iA�T�2`�Ac�WKЈ���|،{$ʩH�<|�����,���e��\� �~6��<�&���4g��0���2GVZ �T��f��NU�Sd�<�QW�"�ZG!�QV�5��Ő�-�h��.�(5�k[Zװ2�m�+j𖾨 k���nna9���Z�n¦歩'�3�萙��'`ze�mG�\'��F"
�6�t&��k}"��ڃ̄a5w�1�M�:� ��;��8�����n|bn�J%�'Sc�J����U�zӿ2%s 8�|ؓ��;���
V�6�6K�腬(]��L�[+B��s8�/��Mo����| �	�(�~�Vt
�(8���g8���T��������e����vWJ%~�?����<����'���)x�D�Tߝ�X�y˔Z�CH3����{���]�Cn^i#1{��D�����O���߫���2W��bT�-��+�ӎ���h���$QfwI��K�c^�~Dz'-~�pI������ɏ�Ѻ0NxZ�h7�<�L+�r_�A'!
!�l�|p�h����n�
�hXmo���,��L��[N���A��<5��1r?�}��u��&0�Z繦�H��������כ	���I��Q!��!����<�������拔^��u����S�|}����|.3Z��[��U���`�Am�Ϋ�����C���N���ZV>�G1���!�f�t)��ր兩�����c��R?$w��=L}n͋�k��6��ѵ�_mN9���G$i�3mkXP[��

�uS�f(q���eJ�uina���	/��%��>E�S6W���	���QTǃ�~T)ѯ?��\Y�Li�?^�%���h���76�y3D-�Y�l��Oj�?9\�W��ngjqa�L�ࢯI�����f�?�����B��"������� {Fxcx[q���b�bSg�|��}��y�5���Q��x�'\��مܦd#�Cӯ�D���#g.�,ۺ�_g�wy�O��jU]�k�LI>Y����2:w&�+C8ŋ|w��-z�ߓ�>Wv�X)�:��t��:�ѵ�l��[�)\`9�c+4�V�k�9ѷd����)臆@L�9h,Cňy�٫o
�]�����p�ᓚYml�U��f�W)��+V2m��T�cuo���ZK-��F��F~�Xf��:������7���ve�*m����jo�E��vp�½Z�&�W:x��1�<��9@���Yr��XH؅	*t4wB�N۫{��J�IN�5�)� ���rͱP��e��.�M,�h�
!NW�he'%N���fƊvy�^Gj�v��qC2,��C>��U',dUQ�~��By�Rں�qb��7W�>>��s=w2�&:QY��`X`Q�y9j{�z<�u�$�נ5��O(�4�,���%�^��A���������{)�\�Q�*���d�[��W�{��jcVI�6��C8τ��`�fX;,�L�ĔS�I~2����m<�r8�i [�4�FflX(��Y	um�[�o�RћJ�Q��@�����]���n\F:> �4���1�Z���"^9��h��:
.�4H�(��0��u]aَ�x�e�,�E�Z��|&C"��^}��Ġ��u&P�ۖ'��VKB�RU2��
NKM[E��/A��u�]{b
8qm�jq�&�H�Z0�L��=�!(��&�YG������Wǚ��h	p2K�Pv�jN0#�'d�$L�'�R%��K�h5c �����8�����A�]\�[����൚� u�E�8��E��jj"w?�#�'/�� "����?����-����~u�������r�7f�|:�����\��4%��є�ɯ(+5��FFb���&K>�6̿w!�_�Q�&���l�v��yb�dmS!��j\��� �[�%�7�"2X8�P��a���H:ؚ��Kkc�јD��S"�
�x�w���+CS�>����룚eh�&���h�����%��ӂG�C�|�� �&LN8��e�\S���vs�3,���m�h���2�G,���-*��JSZ~�/t�k<L�Q8r����gΔf��U#�t��6/2�h�_a���x�؅Mw_e�hSN̙ǐȋ�$�@-�rS�2a�Fꌵ��	1dj1�%7	Z�+��~2���9�����˛�~����@q�oK3X����,r�J�-]�{�]���D�ʶq�f��G��:-B!�X�����.����4U��m�h� ���	�P�@�d54�tM�q�<�,V*�<�a����x�}�R�h�L{y�E��eڊ &$��<�M�b�gH��?�ȿzY�;g:� m�LE`?��*�9��EQX�l���e�d����d��P����>'Ƈ��*}w|�kD�/�B�����5�vUMm<�º��j��	*Z��F���?�!9���3�R^�e��V��1������sDwO�����z/�xo�s�ɂ�D�2p[p{7�<����(lԗ�n���:4y��&gf��A���y$'i��qBq�ݥ���d�r�ڼ���Gm*� .�َ��.�JV%O����O�����ׂ�O��J2caK��Z`�$�l�P�'.|���c>)�?��$)�-I�b��9�Q�8�&1&����_z��h�|*�D}�n2>|�� J�ƿ������㾒�g3p¡�ڍ[�"t&�/>�13�w`/��Qv��G<si^B{��P>M������Շ�$x2PU��t��áO^Xz�ؔ�C���r*2���c�Z>��O ��`Ԅ��e�Hh�K�8�Q%���^4�.�]�UJ�af�@�o�ℏhkScdw 2g��K�1!EW��]��g Zme�v�!>�X��Ļc��]0�V�������g��I�ُ�<=�h�vjhrqE��6����$?��!oa�����eI,�h��z���h�k�/3_A��o�1��y�x(����XV��1%�0��o�z��R���{<i�C7�j�?����2��i��E ĺ]l�9�f�~u���iT�t����`�Jd�f�	ý)Ww7miLjZ}g6�q�Xf	���W�Nx���Qi�o�4N��k�����i%-'y-v:;�d�:5un"G���!��&��ڗx-vc�tk��'�G���9�/xJ��9/��V�l#HY�8�����ۻ�\�c����^���$�+���|$�w@H����6��(w�����C��d���{�y�	,t�� ���Ԅ�LH����ޒ�od,7ͺ���W����j�0a{��rO�:?�3��zZ��!���j�d]��O(�����5�����:a�#-��k�*}�-��x�U�6)9�P�J�-#8���VTu��5�N�5�}��@�q�����+�0+=�b��smI��6���y�%u]�¶Wj���8����I̋g�M��j/�t���	m.C�0�/4�&[RT+�kT�8�l���j�Ǟ��m2�{Al�H�y�i��'��[��eE)�������p��Gcްv�3�j���I����N`�`�?�r�W{Y��셔�u��R�8ܞ��o����K�P,I}�P�!��R���Y���P�t|��S�(��.��|(�S.�`>�AmeRX�t�yeFTPn?mh��� }>:�e��uԠq��[�������^�E���xJ�4&!)ˑ���ʠB�(H�!����Ȍ}�y�<�R3�s<�C1D=�d��[ �*R�5�׷�mg�W�g3�[|�U��(�.���!��<s7g��t�V6q #���RȆ��ܞ
��F�������R�ա�1�)1fNN�b��v�is٘!'��lm͓6;O��J�gʚb�f�@xO�"*�W���.����[����˯h�,������Q?��@��s�>nt%�4��bn��h%A�=d���
��+����usR��߰-��=ɽp��)!X#Ft�!C��g��VzѠ��4�ψ�"4Fp ��3����pxx�K�k7�yܳ�����oj��$��:̵$�w������G��%�h/�4�x6v����K�`�f�O��G��|"��vo��oU"�=x��J�tX�f���܀�U�;zeꄝ�D��o�J���H��9C�i|�i����t�Ԭ�Q�����^V�� ��s������g��?�-�r����.�e����!���^����F/5�?�dH"?ش�T0(�z�Hlѕ|3�d�戶��FD�O.��	��\��
����W��<��d�������Yv�$2�������	^�wG�p���K�Fܥj+N6qɩӚ�J�� �V��^͎-CD�+@��J��}�T�`s�k�v���[��������E��;d�P�,å�!��|��C����;V���&���<a���ч�iC���^r�NǮ1nCO��A��k@�F塅R��*N���p��vg�d� �6���梥ģZ8�����,�*���uA� =w����?s�\Q��jԒ�� %~�׻�R*y��{��hĲ�ѫ��/.�h��h�{��F~�:�G��4Sgx}Z(&C�\��5�D*�~I�l���A/U?(B�Y��uX
/�E+$v�Ie����n����ќ�!�~ }�ѿvxT�U�n���<�t.�~�#�U���Yk�N�D��wy�L�~��\�΁��&�}���T�u؎��y��1�g1�5Jءp��A�[밫����5���fذ|��b�y�l0��g������ؤ�^#�B�a��`�^|N�q+���Ү��!#�e�Z�lg2���.Ҝ�`VR���5����T��LT�	��s$n\G�*���N{Nӕ���ľ��^�s�l�8�dO��yJ�����)�@%��2.��<b�wK�]6�G��T�����wH��3@�\�dU�/bo�[@x����ö� T��a�bq�{�	V�Qz��҂�S@r�~��W������+9Fk��.7�`�6����T� C^IN���ٺ�lf|F'�4�*ލ�a�#95�\���U��+?�ζ冮��&��68����5 �&t{.-\j��Q{������c(d��:�K_�� �Td�� ��a~�#AUXI�`�Es��'"֩9f�pTq3Ɣ螎S-��ۏ�0&��0`ys'��4�`��A#��p+fI�0\t�/=i��=����a��,�5>�:�/����Ԁ𙷑<�}I�R��6�Y���l%��T�J��Hr��|GAe�t�i���:C����"�܆^t�C��T4�H8/��23M$��2}lt{}���� d�]��������Lg X�H�h������CZ�8h	4�KV�X�}ٲ^���!�å��1�
d��y3B�{mfXS���5�qp�s�t��PU=�����x�4�.M��SK)��BZ��dEI����8H:����ټ�Ǳ��rC�ڢ�����b\6� �<���Sq���[����ƃk}'h�f��5W�� P�<��E� S���pͅ�����<�w��Iv!Qf��O��@��^�6?���V皿�;Q�F��۝���t?�I�0�Vt��P�'.�l�W��~G�"������r�S3�1c�̩�8�,T���j���i�?QP��k��p�;6TvQ�D���X��+Ǚb������`��j��R�N�%w @`�}�ϟ�qv)/�^�SV�,�X���=��t���:9��<�\3îfa-sC>z��Y��l�e�"�ڒ�421��H#����ڀ���jZ%d�r#(�O�$��^��d��8WD��g"�:�'-�q�ĕ�xi|4��.�W��R�D\�jL5>r��}�G�s��m�g��dӛM4�/��l�yQ��@/ft�!�{%�ہ|��Ow�#��q����xi<�o��E
��(,-��ၓA*�q�F�nu��'��\?�B��Q�袃o�mΙ���u�O�B�?�@߳�����E�~JZ�k�j��01h��>6�.X����繠��� ��?�;7 �~Zd� �!�r�7ne���6����˅��-Ҥi��B\�gǱziN�������2����6�v��Ւ!�>��?Z#��U�55��R��s�>���q�H�A����4,l��#STY͆�(h�6��J>�\�Ɔ?�t�|=��N�u0��ce��'���oVx��dRb��x)�r,��>Ի�yT����Kt� �M��p.�i�eF�dE��|��O:�`a�����HAzqN�N�������p�P���u˹t���6Z��zd� �bU{	���}χ��=iB�Nh���.#'�hn� �$�]$U?w��$F�iZ���P�E2��H/{=(��J�nzp��tߢ��[p��Mȍ(��-9���LP�?���~�4�U���$���!�jN}i� Ē��^�T|U��!FUz�.@�*��Q<cw�|)�0�����Hn�T��Qx��w�?ީ$ C�(@�u9�ħ�n�UY4�|�żGQ�m[z�a2ZzKD���
�jw!�-���0�4Y�~=g�-����խ��~	��U��A�S�3P���Ǚ������G�NzBi�l "<7��	p�8�/�>�Z������i�uq�P"�+�1�����
���!3ݞ����9'n�OQ��IjBzx��̪}I�E�;
!��os#afK9E>�xb�����$m��[�ǐY�S��[���!�qǲ0�u�g��v0�n��hw|�t��\�2ΐ�SP�қ/=KD����;�i�l��@�[#����m3�':O��p�`�-U�ی>xjLf��@a�>Rh����nmR-X��JHv��c %V�/�l���2pg�y�p����Bo��\�kv�P< ̓�������B�	䊫 اq���`xT����ͷ�~ڷ?&>��1��Qu�@�)��;���F,7{��C���_N�3O�z�d�xWM�f���^;����e��d��Hb����M�Iݺ�ʖ�������O��7Ġo��C��V�C�N�T���J$E�
��$���:�効����Ԭ����X-���c��A$��݋���
Ekie�(Gj����|��nLu�<DopXYy�;�&�U����-ؙu�l��??���}���r`�<1���4�j���_G����-�c!#4DF*_ފ06� ���#Z˓�f��f��Qy�2��ҡ�M��B�Ѱ<w(�]�_�r�E	��=�I��J �cZ�"j{�s��xy��6$1>���	�E�{xjm��lP�΢C��1/�&�8Z��A�ǴO�2��b"/�8	z����I��0Q�l�p�:a1�"7��kG��޾���OǷ�Ѽ�=Y'WH����Hp���'�צT,w�����	d�u�H釃��ё��z��c�M��(����Y\g&�݊��]�7�{>��p�-F��݀ޢx��htx��)�� ~��ô�$
��e��u-��'���Z�wJ��,<ލbN�e]Ы%%��U1��Pm?e0c����9қl�{�X�택�q}���Q�s)�\��&Fl�u��Yw?nZF|�m̅�G���� ��/� �O����ޕ����YXj[k[U�+p�Ԑ�1=^�kc�H��A@{���ӎ9�{�]�- d��/T�1/�U��h�@+�ߣƺ���Y��y.~��4�8�����^�7�4��tV7�-'�}š����&�:/*$���걌5ܪ-8Xg��b:������wi`������t?M���1`4'!	TB��u�:$���(�׏T�`Z �����t��F��vD�7��`�q*كZ�g���٤�&���r��:`h���6o���P�Pi�BQ�|�U2�h�U�C ,����}<\�H1��+�E䭉zKo�0Q��s��l�Ev��a�Q�6Q��K��m��(f6�x��>�:"���8E�T��o7#u�B�&7��K�(��K�]0j�\Po��A�ގkx����j�x|��X�^1�)�tN8�J��D]�q��oE�Si�&��X�,&�z�凑��V>��%�sG��)�zy���Qy���:�Ou'<[p��H�F����@R�����l=�q�}�u�ء�(���K�G� �x;ˈ�Ŀgw��k�Շ8�mr{��౟����bi,��I7���?v��E��������!i=�?PċQ�7ӊ{�;	i1ME�t���f����)�r���y�vئO��^u��ma�i���V�*�k���z[����r������	y�yc��u]��V3O��.�+�k�@�]��\)�'�S�'V%6�@ʇȢ}�k|X��5\zɥC�T�5��@��K �>��w�-C�3�K�sl�Ч��%�S�}he�ܯ�T�l!�'}�*��F?�9bW�k&�ۣ�k/=�R���_=m^&�.��G�#R���m	_�r�x��#��5u��;.� �Pi����',��DVI����N�,����kGLmh.ގt�|��X���I9$C�	B��^C)�8`TƦ2�,����߆Rl���U�p�v.�j=T<�ք��KXK�-VF��Z�Q����1�'~G�(����%�|��3�Q�ۛML�1�?��ɤ��xvVq�  �Ϧ��uZ%��g��6H���� ]�E^�*�9��tk��P������h��f�[T<�f�V&���k[�뚪�����P��v	|���ʵѕM�5����T.�՝{�$���&�n��D�+��i	�m(Ю Y���ʆ�|��?J��C��7����h���w�PRU�Pu�_8�Gm�~�*�#8b��,��ı��6w(2��5V�r���&�6����#��n�.�\�����������OC7<��\U���"I��L��Y�a�y�6!5��Y�
.Օ��дS��^�'�bg�:
��4#����Rs�?,h���3�@+�e��
�q��X��u��V#$�*��2����#'��"u�I	�YZ9�U�u��]y*9�����BQ/����j��emR�114�/�	]�5h���SfS=O6�����{�P_W�%iM�j�0q\\R����S�}ਆ
�a����3�Zm�8�$��$+Wj��̨����]����Y��K���}^���<�3���Γj��>��t�5v�BD���_Ze����K����;r��W3���!���\Eړ���l���еN�t���������(���UTq��ȭ�Ij|l�/H�=Ʒ�:�R^����wwλ���W
F�N��..�FoR\K�U*G�����=y�e�r&.[s�:�^r�q���e�9|����Χ�����������;N_f�n�q��\��l��������r<W��H��DS��-�|�v?I8����0q3��4Z�3r�W�(�3��QؿRӛ�N����]���˱��ޟБ�I4yV\���H�@D5��*�˶pF���.�K��L�鸜l<��lL!j�����`Ƞ����	���/Y���|�'@��@��V}Y�Y��28��^.މw'��e�C����T�Uzxk��Q0J����̵�@q��zU��ICǯy�.�
����4a'8�#m
d>\���l��O�ddȈ^+M��9R;���dR���/�.����T7�-�X��r��_� ��� 	7^=&×�����U&&����s�5�l��ٺ��.%��"e�+�'���0�^�6 -��=����ȗM|Q͏���z'�v���3���-2���B����_!�Ńk�Zh�����25;�db�R��|p]^lM�Vj"�{̀�N��V�%@:��`��iI�u�dB�h�6@�ЗAi�ЫD���`VrBt���.�`r*��1��)�mc>���*��a��A�;���^���W+Nʐ�����V��wQ�H[�="x���B'q��б�|��JYǪ�4yʱ�y�,����O1.=�y�ս��A�w ��$t�a�H�#���A�ב%J�m_��Hu�>�:��S�/��ѷ��̌n>QJ���؂k�r���-(TCk�
����&�	R��<��G��n��г4�r5���Uu!vAn�	T�K�� X�<$`0�.�gWԘ��s��,ԇG�o�ݬ�%�0S���3����&�W����yq��H�ߧ,带�d����J1.�3}�+���<�m,��CI5���H��ojao�(�N�SvТ"QNYI����7K�Z"JRP.�H��{�{*}��2���NR�Q�
��ޑ��a�"YZy-"��Jg3ԁ2�(�色o\�G����|Jy�w"v����$9���3L�>|���Ã����3�M��.-�o��Y���{�cJ0��[=?�3�˙�����ؿw���\q)s�V
�����\<U��� �!a��Ғ�9�S�k��q�k�]���	���7)\%VPH�Q8~
� ��*��U��{[�_�8��S~>�l?F��l�^.�g�`��[3+�����G�J�Ӗ.QO*��u��!�^������G�ĸ�mˍ��v�}�M�u�%e�.�lS
ig���M��H
�u��H�����e�Oݚ���+�d5ۋ6OK��؋j�)ϫ��d��RH�L�
J�,�5,���r.��eRZ%�R�ې*�����Ax��9����'�����A����t�tV$��r7BdҘ������&%@�`ߋس�DϮ�D�Y)c�xI���J{�?7��ɋ])5ag�����C7 ���i�K����­�Ȓ���g��4d���
�����9���L�a��n�T`�K`~|���J�_�6�_���Ou>�\;�ro���Br�%�Z}�:x�-��P3�6��]�[I(�$Q%�����v�}7��GW:v@��7��W���)�s&�PJP�a#���>��+-,@�m�O����o��.-�9l�@ةQ�7����hv&���kE�����Ir��a	ǎS/K,A��Ӥ��L�
B���3�:3�YmI��g5m'E�.��#I�Y������\/�C4��Ѭ^�D�b�vm��+$/�?'��Y���u��$�m���x�6*h�+�ʎ�(�����W'�'[�N�uu�St�}����E�u�'�8�sd�`�U؛Q�Z�<�zg�:/IL_U�qK���ؓ�4B/��|i
�`�KX^���hՒ OR�#��D��gZv'��J��̹�?��|s~խ�V�acፌ�S.����pө^�>$,o� a����֤
|�>�[}L
/�,��(���h�W�!erU��Ɲ^E�+��W�Uz�=QkI ��r:o���g�q���������D�����fơt?^���ڱ#ᰜ�F���ؾxTC����o��z�/�^����"(MbB棘Q��z���ш:���ji�İ�u&�@��%7�ZD�Y�W�[�h�5��L�U�ٖ^gQ���a��JL�e��;D#l��g��ݦ�c�M��9����p ϋ��S,�,Y��>N����ͷS��ʪr��@\p3Й��¹�4�/����x߉�X�]��z�x�7�M�|�SSPȄӽ�q���Fd�l�.�%�s;i�C�"��)��x�Nb1��w�G� �8}�U�$�h�А�Kg�F+���ۀ�\��%�%KP���IMl��sOvXI��n4Ж�PO�8�X��h����:#b���>��t���ȉ���� }���U\��&�{e:���w<�hu�@ڒ�9���.����N�1���F��	�cn���)��oJ4/[c��U�k�.�U,�
�>΅}�M���
x��� k�qr�!:|&��w�h�PY$���>7��{O���F���?������Oxjx/�����"�7�%w��R����������	 ����( ���5:�^d]��W2������Cew�Ee��AxZ��(�M��jX|�p����P�V l��e���4o.4e�y֊�@��>����^�Q�|#pо&w���գ ����FÛ��m3-�f���T᮲��~�OqS���ne�z\F������ �>L$�_��~jx��JѺ�$��:�s��p������f/�/C��*�x��G�O�����d�Ǜc�m/ 1*�9	G�����FF��m�z@�,!��(y"��r'[9��7�����аY��p!�3�$��lU�Q�1PI����~�Di������k9������;'59���2ڌ�jEi����Ss�0��똯#ud5�ߥ;	$Ǣ��$��	�h2���ڙ"bB/r�0J�_�F8��L���eh؟��Jj��&�QGe�
ᴘ�%^(�0e'��&����քk�}b^[e̍�l�C�ڈM�����'�B�ڍ�:�m�f<��6&Zl��,Q���ڊ��SS���xp��p $''�<$������)���j�Fͷ��w&C,�|�H�ӡM9�HA[4��Q��x<:�;�B���vj�B."&�hJ�v���˨>G��K��LRib�]�K��ٸ�6݅�[� ����x� M�?�p$aT��ӃB�r���� �Oˢ�f��� I"����l�x��N�0�����NC.8����U+���K�WIa�NO���|�f2dzQ�c��W������*���+�.r[(�B�%<�������c$m���A�^f�;������B!��˻Ѽ�����%hZ��}���dL�%]��g1�N���?��3��]*��f�*�*�&A����+	�Q�i��������DBN�}[�0��_[�r3�*O�Ӛۆ#sHc%W!�g���aK��9��z�+��1$��ዊX���&|X���\�r�Ӏk��u&���5U���z�6#Œǌ�_�`�G�ۑ�Z��~o.GK�NoL%'"mc�
��U����$���[�<�8׆8wh�$��P��N��+�ӧ^�2���9�9�&�郺tEg�74ъg�W[Y&�q���>����y��GwҤ���0Lʩ����+�OB�U�;�*`c�&�z}�dU�W���&�J�!��.�Ә�Q2�Q%^i��gڞR\B7�+B���n�:��]7�[��|2.�0�g�s�@�(�u���-����O����y�Z�|�mϜM�gT�_uZd�l+V�-X�#�qT��H���t~n:���Y��6`La1��X+���E����m�� ��@3����j���S����&/��M7��橥�hg�O�X�0	e\�0�P�x2�#�r��/p������Y���'�]�9���Ыቄ��h�/���h��O�$c�XnQ�^�Qf��ALsR=�%:}_��&��O���}~ﵨ�:� HV��@K��c���i�[�׻���S����R��~/�a	���3�.�|��^#�<��;7(���]g�?R��SI��s����pp;���?�y�t��+�<����'�6W�Sܟp��*0�-wi}�&p ����#_�G(��/��FM�������R���R�
	l7�)N��rx��>K���>1�)-�fah�/,zyf%�
�@�^:�2�QeB��X<�;���a���	.7��j�:"8��JA��Y�ރ �� Ò�K�c�����B���Q,_	Qn_Kפ�)���q�8H��꫃ޗ���)�� �J�b��P�J��A0S0�/7�|pvH��qB*�Ы�J���`�C��5��V�Isp���z=����5��r��H�L��'���:�c��٢Q�k-"���z?˩�hh�0���.�M��T9 ��Ŏ�`oF�H3-��U��	���fq�ǀ���]��+��#�r�ޛ�Xd�g�K-���Z0<c��5(`{�!��J٧W�����fF<��<m�I��b�'�n����p<qI�İ���5�t��┈�p@���1��?��$x ��;�w��U�"�bj��#�Vג�i2I���M�~�N/�"��������J�fT"�a5f��o����6N�;��)}���1�8�������d}PLK}#�z��0_y��|W�RK�w�����x�� _�Qe��k�q�v�v[р�g9P�<r4��k�$��ھk����q��[�q z������R����#Y���n�)�+0��C�kZ1�n$�"��n�G�����b�ފe�/�f��Xٿ�]'������)��E��ĸ�v�<��jb ��^���	��"&&�ؕ��j7o�}�L�c���X��z�8��\���[s#�&]ўNFV�*l2��a���>yV�e����H�it�z�l
��R朙_Hv:�2cp��M�v����Pսs���K���?[�Ls�=NK����B9��m\��Ra���4p����A�|��쉄�(,_-�G?nҬ�}h<�j��×��y����m���`����L��j������(o�	�=ICBS�Hs�@&}AX�rf�u�����M�P����_���v�Qvi�XH�E�&��M!	Gcr�Gc�n��s�q��%�t�A�u�#x�TB��5f6'V�yˮӿ��}s@�c
����db����\�4^�r"\C�5I#�#���j���@������1���Y�ݛa���>R`���źx��lT�{�<%�+�p�`�*��W5��.��Q��x�9��Bb�K�:�*x5h��N�V��,�9�d,�w�]2�e�c������m�����gLT?s��6!��w����Xʍ�ɦ��(��%`��%���!ݣU~]\��I�E�|Y�$F��\�d���9k���ĽK��ҵ�[{�ao1%�zY+���a�x����e �����C+�ѽ�{�7�����gT=r�i8����g���dR�?\
�(�TF�<��ۇ��
�6o�e��¥{
V�L"��t��\���خ��=����!��U�V�1��9a����8�Z�P�KhG_�����z]PR�+�AF'4�cI"0H B�aO� 6���������6x� �톿k��p
<���C��yJO�@T��E����������64�G�����@����"@�q�N�S�o��b��O�j�m����2n���稒 /�CL{d�,��{$������r�.���1o�h����fH�G�c(.��F�;̪*A ��qr�|�������,�(�_�������[�1ԩ����O���驑U�E�+���o{� ���'���}ۘ����� _;�V&y���n����k�hG��!���,�ޓ��#��\`��'yH^��/p�Xz�h��R�B� H�r�f!j�@�ޏM!Ƨ�ST�.��뻑�{�����$m���Z(�π�7{�W�}7�+�Q'ף%3�U�F�bt��0����� �nӱ����t�&7����ѹ�Vep���u��:%�)��8.�#k<%_�Nڍe.���8�o������t6�+�y�ԘR-��i�+e�@J]��x�=�z��_�'WV��{����<���G-����̕�d�cg��?g��6�7(���qG<dU[��<ʮ[&�Oerå*�Cy�J���8���EeC@��gG��+�$���t����|pk����T���S+	k_[긳�ߝ��N$���()kj���[�7���O9��/O�p)�S � �G�o�ʣ$#v�����<ׇ�F�?��a.��=���x5�[��j�:嘨�3�5�S{�It�q��E���hնE*���`�V)�����sP��� ̿4��6ZRw���kv�rZd�i���kP)��L��m@c�A!��;�
���p^����ۂ܌x��9cN=a�羵\>�Z�>�5<pdR
�k�LZ�$s��?9ҙuX4�w�g�Y�j���C�B��A��Wq+E~����d6�lFR��f_,��IKf�B�����;ӌ�t�J�/�˽�x��ҧ��ӡW�r��͹�.��>?>��T�kv�4h�0�H7aQZ��	�O��|�F@|��/�R�%��Z��ۚu}g����:��J���� ܻŴMv,Kl~]W!�E�GK�Q��P��^���qemh�X4�^~�ػ�Y�z�G�����5d�OvlB�h��2U���I�,��{23�!&�/�a�����w�BU������&
�}J.y�t����3�&��s�� pU����!5(�{�����"p���Ή�׹�@�� �� ����M˅�>{�p�^����7J g ������n�I���y4bLf�+�-����/E��)(s��d�{r ��-��(�˘&�ޮ��˂�@�*c�d��x:>��$�2D�@��"O��R�W���Ft]b8P��Ӎ�Ɇlr���ˀ�n=��E���:�7/cl��V���c����0��쐭l{��Vk��JM�?�:#��;K��u���N��!k	iHj�
`�f�2��k�u�qփ�z�a���}�̛�X�@"1���5����b6�|������>%(J�����cX���j��םC"X��,��H�Q��6#���RG�"ŭ搦D�8R^h��<�*��b����T��%oB������;�����XLS����4�ƀ�a�S/Q��$��#b~�	p�=�=雪.��� }�`�WN=��>����n�`�Ƽ��]* ) �ʸ8�yU�0��v�Fm/�F�3 �q�^N��q����s`��>��x��\�� ���N���6��i*��_h��>n� �C'W���[������ <D�����0��3����ѷ3Q�=gg^���]�R��Q����
�w�;�K��.�L�N��ڻ���pE�I�4�(i��?�g`�\��IܨB8,�L�w��+��*�p�#PX��Ȓ�&O ��iŅ�~X��x�1 �Yj��0���X���"n�F�ɩ��j�Q>�湒hM��5�Z��D��%�+Z���=���znT)��O��U<3oMV�r�g_^{��P��~*�06�v������6|����%\��8�]Y���[Z�3�Nm2@ca0[�ʲ��'�������<�T���]iz�i�Bl9>� j�E��؂��50ĝ�Յ�+ܶ��@�o��r	�#�I�a3�S~A6����jT�O�ⷍ]���,۷M([� z��<�Λ ��$c��|�A�N�8#�o�W����+H;���e�.���`-�Z�q�@
�$́��FM��ؚ��te��}E���Q���n�A����e���`S�� E[�;�u� >�ip����"X�JYJ�=+-=곞G����X���;�H�/�B�S�~�dQ�EhpK��Az���>��&�j�ǫ��	Qu�F<�����$�>`U���S���)	>nQ��-"XAS�V1�⛙&�̙#Uq������#�z���<	ǧ��#��+X(�~ۇgZ?�f}�<���~���\-��9q��>I�m�WY���x�t��K��}�����q��y�&+�Pv����Lf"_�7S[��B�� A���E)Ѩ�j� �i���a+ ����3�=�"g�@�Ү�$%�g8�`ZJ���P3={B�T�n(|�ҽ�ΝݷZF���t�����Mc�YB� ڛ"W9E������{?���%�e�I��8@Li���qtO��wЪySfnґ1�ʂ1�l�o-$�\�˵p��*Spǀ��#�cM��i5��=�̬��M�J&���A��I�f8�E�xݧ���s��@_o�!EC������0� �f?�L��13��v���%twbb�����ݭ��� ^����!؄��6˻h����b�(�����=.��o����w����n�I��H^瞝���e|8ַ_�Z�?!��!���v�Ҧt#ZA��6	�Cc�B�~���y��|�+MڰF�(w�� ���<a��B���L�m-h��8@�qcct�ӕ#Y��L�T��o �Q���	���?ǅ���;���+e�h�y ��SCO֔���U�i^�5MDש��M�ԖUh��a%=��Cû�����s�
:L`"� s7��qN���1���\x�y�V����v ����/�#�)'�'��n������# �H��cf8^�\�aP�#Y��NzAw��TXv�oÄȘ+�������~�8�Xu���:ܳ	%��AU���$�"�g)'�7;�;&�~�k8E����E|��A�)��~�UI��;�N��}(�tH��3$�|o�(�t�����0�2��|�4�i��ƑfB�F�u��|╏Zf��r���/��n0n44����xh����}�RaB1�����@�q�+���p;!;3�m�ʜ5����u��af@�>��CPw�z��bd�\$�#�����V���[��i������cT+�9���;�kih_\rr�!=:��\J
���N�ɸw�o�ӶOk&�%-�-��"n���r*������Z��4��q���2�7�#�2���Bf����[�5*Wq���$`k�3I*s|l�4��t�O��5�Pv�تF�A-L�f��pB�`@��.e���Õ�n�:$��_gӦϻC��t�:$a��������{[Cxg(��j��8qP��z�q�ms�|T��$k�7�"�]�����oZ��+�eH;�QIaۛ�����>tz�E�y՝-�}r|�+��+��<��d���YG����+��ь�r�],=n�m�P�n�t޸BPl1|�>	�8�U��Unӷ�R6<�:|��]T�b�d&����qٴ�n�&�q��ؘ�V��H�?F�c��!�țUpXuXx{d{�#E
�o9r��`�S==�����8�����)�}�4��lp�Wd��dC'�O�D��@����@��²}�0^3�WO
�)�f� ��z��(��Ha�"D)���X��8�@U��=�?nS5�������n]F(��	�������ޒÍ9�g�C�K�I:=��]�/�~/A���]�m�L89�-��Y��W�:��m�&5V��i\)�/�\�h�#����b��/QUz6�9�4c�r|���Մ��Gn�����w�-x���ǽ��h�m��p��B]����7ԏ��Az�P��t-V��+슅%<�Dn�p��Uf��?=c-f����|mT���g�E?�vR��G���UG��S��!^U׋��$�\����[�=H��q�O���� �v2"�w�IVpD3��"wݢ�/^V�I[�t�|�D�V��ꇧ�R��G�����Ūf���f��j�X�(yΙ���<��O��5���p�5z�ǧ�{�*_�0�����*1�OH��?���VH;awM��I�o}a�Ǎ��}/�ɿB�����%�&�x���CŬ��9�()smݕ�tU$N��"3�ř��3�Ң[�������zAHh)��K����~@��~X�"O��(�O)p�.�yQX�d=�Ab�ظ�toG�/�	�2dt �H��dY|�O�Ô+\��0�����,��_��F{:�u��c��̳eC%�NW�eG�D��%�ߔ�������m�ɳb׀�.U�;�,��}�G��S�����\2�j��P�L-!�kѓݔu�FA4��l";���\4$�5�q���;G�w��o�֬p�{�����j�E/�j"��λ����o�]]���S���m>9�>M3z=� �)L�؝M��~[~�����!w��U�f�7���
���	r����*������h��z��ϻ�-����9v�}^�>�(���t����U](�'���8�k���<��� �&���^gA�zK�@}m�dæ
u�M��-��Ǹ��Y�o�t\dh�4�C[��c��d������h��L��n������@��{
����6ٳ��<���*����M�C�.ѧ��2���UL%���S��M9�+"UUPR�´�dX�K��-��Y�򅀫(�}��R*�6Cۏ��Yf\�F�/M�Z�W�E�R2��۞��d���cxrѐ�2̮�K�Z�'���1,�QZk5��Yߚ���eu�4��<Y��Rl�y�дj��q��9��WRv���[؝���u��=}�-l\���"��)�n�8�B��,�Z2�����\�nv�h�Ù�Uh�4���8���l��S���A6)�N�*��|�ɹ��e�� ,�fz/���'�A�`]��A����im[�WݦBg���]%������^��a�W.��cr^-RA<S���*�"���kU�~��/c:�A�)@�h���e#�㊀Bf�=scVf&��u�v���j:��*�R..�HI����"qE��[�׻���b�::�����p�]���c=���;���w;��6a�f"�	Ȭ�F(T���I+p1� s���X�Pφh�EP���L��?�C�L��s�����MY��ګ��u
h�}]�	�%{�����n���D�!��?���j�1N�m-p�m�Q�Td
�a��~�!o�@�I<"n�4G6�fK���L��ݾ��Z��HvG	|+٩����5F?� >��ė�k�P�
09O_Hp6`�0OΤ��o�+���U�J@zQk��*9�#����G�\, �垩�29)�4�Q�kd�k�͹�����)��ʩ�.V��x�/�ш�w�����w>����>����9�5P稞6�#ZL/�i:���l� ��&W	��U�ZF��kݝ=l��tņQ5.�g��8�U���;�ߓ����!֯˯�`&y��E��=�kKP)�rú=�8�
_�v�^�Rv(Jh�����|��Y++9�Vٹd0(^�N�8id��-=�%8�����T�Ƴ֊I��G0;Ѧ�
e}.�i�E�������k�ip���u���<V��a-��*���,��ŕ��	g�^MR-�0�o[ =wb��Y�h�Q��9���L}2��*� ���{�� ���*/��9v�� B�nV��|I�țL�Gc��c�������*��H�����F8�앃�ʓ	��)i�u���A�(k��^ʕ9ѩv�R��jǌ��lx�M�?W�Iw�#��J�䏐<���{2@�Y,� l��g�����f����n5Й����H�
���U��\N{�<*w��ӿІe����)y�U���M~��t��|�VI1J^L1,�:̛H���Չu"%�H�oWN����n����&��@G*��ش�bH�"�@ܕ��X����E'�=���.����.w+���SX�v^�|7%��X'q)�Ǟ3��@�E*.�]Ni�ً�x��rܺM�E�(��ɹ�(���	��R>5��n$�W8�~/�<�x���	�X�3�P٩�O���vn�����?������1�en��-�]U���l���e+����=�4�������z�'��ȒV  �X�ȅ엂ӱ,�Q�	��p���ǅ.1I؍��?�_�k���\"籠�
j�Yg���ʰ݅0�Q[hM���D��3@'��x��Ō��d�e�	yw���|�E�Q�0��R�4���p��#�J�V�'MA���{��E�f��g��(��_hyS�������G��Y�w�es��<i"�K�,�;��|M��h�yK�~�Ra�*C3}��!;߲�.�C�b�?�Mx���0�wN�o����[:q� 
�_@`s��C;�b,HZk-x%aT�b�I��"(;��Ye�Z�%�J���6�V��8VT�7𷞲����Dj�#�1�@U��ِ�Z��������"m��
ںҬ�Oi3*QL��w����`��k�W�xʦQ�����mf�
 >i���������K����G�(g�&�~�����Rɝ�N��A��v7C{������lH��]#�����:dz� ��D<�a�L���ѡ
e�[��b��h�)hƻg4�&%�{�OƯ�Z�/�;�|��H�c�̸|r��h�T�OʜEh�.N`n�c��qdQRv��F��E��T��SL�ؠ��C�GjR�q��x�Wc��Ě?$���(��l@����ԟ����:5mo��!T�oٺ���XQ�;5�>y ���=����9��,|�58I7�Wg��[y�#�JӴR�e�W��o�~)c]����Ӹ�;*z&�h���}F{
�p�3�m��u�.כ�)�u�O�E����LMt
۽��N���um�Ꮢ��<��/�C�����sV��6D��h��z�/�,θN��9����=x ��w�id'̈���G�>�,J�?�q�A��8�cm�g�^�����}��Q,�ìb�Џ5<RG�{��;�����P@V^IN4�5�YH+����{�É�.K����u>I����f�W���$�9G�5�݃�
���i��S�Q����!�O��y:2�(Ij�h�Z�t4_j~_
ff��k�_Cȷ�pW�DM�>�`�����\�����P�2�X�곻m���4;�`p�F�N�l���wlDD�s?�;�.6k�`'?�L��=~!�s��΍����q��:a��̰�A}�7��qx˗F`~�m�j����B^zcL�o���B��k�p��?�蕿a�0��zרۀ�`h_Q<����6�6�Rz�� i��[g
�U��kZ���ŝs��Q��ٔ�N���������Ü0�[&<I��p4
�2!���E�Hr~L)��V\Bn�\ �f��g	���_o��ҙ�.#��g�����Dϔ��,91rͅ/}B0r@[�]|��C���ZP�'g���B�����L�s.*�_��C���-Q���4�4wwE:�A5le����1'�7+�,��M����0���,A�*^Z9 ���ŕ�5��Y��;�d��ڪ��$��>I_)�۱KH+w�Q^�|!Y,��Kf�X6��H�f`�@	��Ʀt:�g
���]W�Z�m����k�_n�?2)�٫?��%�t���[غ��	�/w�:|�1�ņ��:��l��Nj�4�$��n���G3x��lO��-8�����i�"('%tɸ#A�����4�폔�n>�ӂ�S��O����/�g��a��9^�5}Z���,�RM/&g�֯�������d4���?���S��k�\f�
*�a�M3Y��7ť�Px��]��V�q���_������Gx(�`���&�����S_��O_��,���Ơ��{���w̸���r���󆲻���[�BD�u�����6|��$$5���NJf�B]eET��n^� �4O W�<	�K������|*�m��3�7��D��ó7v'��g�T2q��v�~�ߟe�:�D.?�Lk{�+On���8�{��rn(c��z�t��ؠ,��Ȉ�`�1�Bg4�&fM�͙�d@��]����Ѧ�^j9봢GX��7=��;,�N��߽ƈ;�����I˾�@"#�{X Q'pw�vIq��t���g�ரe����]r�����q�6"����?n��h�f��v;��
"�,*/�2k�Ƣ�GP����a���3AT����78�DF �P�{�<��]��,�p�5�O%��RW�څV4���0D1p%zzM����S�����daK�C>!M"�R����zk/�X����z���I-'�Q̠���qZ\rW=Kî�+�-�v[C�)��Zw� �u����%-���N�H
 a/C�CQ`=]��a��ˋ�T���R��5^�>���3��1���E/�j7���]h�ʏ��c�i.���Ԏ�#�N[�ll�̊.3+@)ӋC�$�ôR��B����n[��?oa���9�ю��Tr:���>?g���?�����!�{�&����!ڛ�N8Yj��&{��Q1��-��_�K�_��;��&�_�QW8�9�Z�`âB��JxYx�]f�-��J���J�,�(��p:�nى�[��a���FrS�?��%�	U�6���e��}�l�6�PP�Y�se�l�����T�ߑ���Y��+�B]E������8�͹U~�GV$�Qڙֶp����?�z��8��w�y�O��@g6����0��;��A�6x
Ȣ���f�mׄ$p3��_� CW*F�<V8��"�d��aV^����%m��|������7đ������|���7��l��h-�â|��ݷMZ ��WrAsL���;����'E�����i1{�`�&��Q:i%��$s�8W����O�vxx*�e����v��m�KK�$��cf��j��qe�D�68��ў����4�yķ�.X
�x\�-��5��:�~Z����!�KĴ�;�]}+���	JMq�[G��kQ#ui������w�+~R��F_��� Q"S8o ��v�9E�(��Z�ß�{�yb:���%{mq���BX��ߔ��B�cD�Xxw���[�ۇ�d.0GG:o���D�d���y���<[��T�_��qY��M=ݪ�૆Q���UĀH7��(��+HT����O>&H��yY�۰P��"��ӏ5��p��sg-��>�|���������A���V�2�w�__#a�V~��]>�	vhsQ�Xo�;�O�e�Q�!Gѧ6�a��jI�8�[�q4N�'=��n�Lٵ.�eJm�f|��*`��.b�+�PI<k$1���>$s�[3��h�s"K��wS��V����FH�M��U�?��p���O��mG	��ͭhd�!s����qq �=�o�Ҥ�_S@V�����"^���x(r�a�kp,�ؖ�XO� F����c�>���E�t�^��
|K��z�[���է ��5�FH]�)s9��"Ӳ�-�Ѵ~N$�D�Mz ���D5��S���	L�h���`�Mv�V���_����E7�yD��~��6��B-�H�|�BS���4H&h3�F[9o�v���t�7��!-�֦��e$s���t'^��OR�5c���QR�),&�KŒ]���Gp��a�)O�綳��]�*Q&� ���Խ<��8��hK��6��-�ſB�-�L ��5/��m;�U�0�7����qL�_M��'�]hx��@7�/�R���Z·�!�ˊ{�Ӧ0����h�6�vd?"�w��2��W�^�>�NQ�{ؚׯTd�Ν�x:������ۀY�����Ќ�dy��y�#�l�����fB�t�]ƹv����`E@)�/s\/���Y �c���3�bv{�Իn/u\z���c,�=3ˑ����#����${H�0���aK|�d�h�t[JP�3`O�:�� �թ�sa��,Ƿ���������~�m4�տ�ઝ�'�I��X�Y
�!:� !��^��Ӗ�]��Y&��eln�� }�uCw	�A=.����1�6��;���*��۵�v��V�1󱾷��)YA��? kR�	j�z|��5�&_�������ɣ�@m_.$)�./��~$��Xmc�n�"܏޷�^[����=�� ����#󁤪c/+�^1�c�:R�-u
����8�2�#�B��n���<��y���M�ܲū�������:�,a�d9u�b@���#�ڲ_�Z����}� ��%���p`*6N�E��P^ ��}��س�<����{1�
�C{:��q��_���c7fo��f�H+�����[���)��b���<j���������$�M����f�ɓ�4+C�����~;�Ͳ���N��Rl&1%?����zj�!��$E;7�R���*����}]u?�}�}��.�e�ٶ]��#ȡ�=`��А�8Mbz����㝜e26ɡYǉ��#a�ٻ�4�R(��c_������"�⿺<R@���ɷ;/J�Q��a�� ����"xK)U%҂��j 2��K�x$�=�t/�Ek�>�����6B�/OL��
�*�þ��#��^�JZZ�����5V{�Z�%�x�X��wl{�R01+M@T'��,�6$�� $�US��d�̚�9b��x�p1���x ΗK�D���2fC?��]"��rA3��GODSm����a�|�6�t�l_o�B��ּ�A	J��-!J�O�we��������݉�4�G��i�:�8,o�0-�g��
�I��L���HA�rZ[����,r����a]x	x�U-�2���O*�'?��h4n�8U�Ցx���[>W�#��H�# B¤��7�Y���윟�ǯ;X��M�A��`r�����d�g6������/�?{"����p\���bEO)�ܘ;�\�����[�ːBܑ�>J���2��Q�"l+(��0�*w�w�1C��j���*�ι�Q��w��~��.`�r�S�� �k󊬏 �Ϸ->t8|+��q�MlNϊ��Z��-��p���n�`�׀k�L���ԉ=�d'���G�.�e�ir]Φ��"�ss�kc��e�iF���#Tc@VQ��*E���np�����_n�11�b�e��cŇo��%]�b���Gx���e�2�J���E�,��
�<��ٽ�YV�N��Q(��+�Z� �\�]ң*�F���kk(V����f��Ǥϲ�b]d�F�JƊ^z�Lu�xx[wĮ)����T!���n�s���<e/B�]�ZE1�d�F�T��F�_�M��1���.�>���`.J�t��ژMV*�H�]�2���f��4	/�c��|��ַxm#_ �����C��{�*Kz󼣡rx��l/��,; �38h<��tH�mƼ'H�s��w���m���;r�bJ� �q����+tQ�W�hV\�%a�Xɦ��v�"P�X_�
��=k�n���<�Nk��ߜ����q�
�[�%��C?���Xl��!Kw���]�.q�����/��@��W�aܟ!�q�d�P"z����L<��<��S���RO�&�`p� y��(n�Jg���]_{y��s������bW�W���� 6_��/t��U����;#B.xNWr�Q�F(���+����x�����G�uI-ԕFu�9 ���=¶]0'�5�H�]�A��!=�6?JOMYW�lOǴ�KD$�?E����◌r�pmI&���t+�j*	������r���XC1v���LV�o0LVö>�,�8� �dh�����)Μ�g�����FV������S�&��f�,A�/(�D����id��_V/�w�Xsi%Xg-r�x��nZFb9���fF&�����sZ��t2�}�p�Y��`KsZ��gӟ�<��S�@И?3��iY�W��zHJ`���QE>V�tw/�,�V�{/��s�G"6mF� n��b�:</�;�A&%½�{?���V@O��G����8s�i}����Y�4�zUǷ~KY�"[�
l�e��6����7��m�G@s�7w�AA����68�	M�P��b��TƵ�P�ئ��J�Hr4����A�u������/�O��k=�{��\�n�Q)<fx�z�C�eyGq����|��ֹ���������K7��ǴPw�u�9,,�͆�BM�_o�qz�_�f�z��1&j�ɥ�h�A%*��CK+�Jg<J���L���H����~	^O3�Z��grt�ȡ�5<�LSZR<��8�4��m���9Ļ�\�Q�~l�0V�*_B�,�3
����9�e�R�/�[e�[�n���}�7��]Կe�B3c.�#�� ���ͪ}��lvP�����D�:���0�ϙ���ԧx�{�#��.���ie3x7)��ne�1&�E�'��f��{�j)��`e��ma�ee�L�~�z�v��6� ��)`2����_yN��i��#����"xd�WGŮd�+�鳫�=�����U�%�o�&=]d'��)����{
���UP������]��w����^��z���S�������ED���tչ���U*Ğ�6��˱[Bk�x�`w3& J
���ߠ�&k�짣Vxa�p�S�m����Mv�=l���8A���t�Rlq$�Bc��[b�ک��J�D�'�CB.�kq2B(�[��Db��ׁ���-C�s	�ؒ�&�0��=){��Z� ����s����.��a��t�y��X��!�4���;ʫ����>�������I��i��l�ȋ�p��6�kB��������W�ׁѺ�H�8h6H��V��Lv�)��;�Hb���$�ƶ9��3
r?�@����E�N)���`Jl3������j����6�A��|w<�,"�S�����L�J���	 �6�ĺ��1%̧����0;:��.�Y~�3�s-���z��D����;du��kK �`}_���0�X-x�T+��#|yˆ�U��?��ސn��7�+y�[�6	;�6�D��a��<Yl@8����)Y����mشh�������A ��`Z�b�b�s��Q_;	�:_ v8b�;�5=���⭊/⪚���>�V^L3�+���~?�.�M�^ߝ^����zD=cm.�!.����O0�*9�u�$��B4����*�6����:��O%�0���5��@6��I���*������A�Cmk���H�j��ķ����Oln�}�Ƒ�yȢj-���9���J�����oPS�w�_�(��p�T��oYG�D�w`�?���Ε��`�g��H��-���0�ޚ��*�����JЀ� b0�m� r�2�h��\]]�(O���F=(�J����Ⱦ� X��W��ʢ�=P�6 _��X��[�G�@��]h++��	�Y�0Xr?��@���upI��@p��w���# ��A6�)��o���jov���'�v:~�J���vx�0R� ��Բ���;ׇ��B$� ���ا���;�Ҫ�cI�� ��)؄��a�0۵����ZtzS󡡙j}��l��B?3��#�ͩ�ߩ�����KW������EÔj��1΀��2�ͳ�T4 ���|��l��1��ü�w>���8�	/��i�"r�']�D��@�χĸ�O%�����\u�1��B�%p'�g��q؅����>���;���k��|yO�9�,b}�M#�ϩ�t�r�`D>?$��%o�5�	
K��=' ���O��)����g�e�"i�a�Y9��q�Q�u���<,��:��;Hl�?�Q4
袘E���7����P���n�ڪ6�ɽXdB1��x{!�ЫƐ#bj�����V|{O��xʡ�;��׹�Gr5���->�j9�*G���h1o���*X1���D���<p��.�
�~7u%vR�L�S_�:d�=ݬ�J�֡�2�-��b�<YY�Lm��v�]O�	��Y�3��f�U�jx���
��F3��[��d��۪���F�⮟d���j�S���3��ngU��di��b��[�ۤ&ຢʉ�Q�~�,6�����$_��j$J@��Y�Z$����ɮ��Ő�u�G:y�6/�������Έ��2[�^�{"�: oz6��y�W�4P�L.[�@����$\�|?�3HPB��%�I�)=��X��C�V����
����^��U�*�J<"��Ӑc��2�̛�~Q���R�z��y,z% 	X~u�H>0�A:�P���ù�5]4��Z�Đr'�h(���nj�ZQ�<��n7l�C��sy�Bw���0�*��;������51@;���ۨF�E1��?dJE��"Z/N�R��4�E �R@��eq^0`������竐Hbݛ��0�ˍl}����x���كQ�K|]=�]��tE���%��f�>H��vm헩�p֜gb�;�?�^;ޝ��d��ܺ3�&A��aVhy�ʗ=�شui�~�M3��F,����r��0(ֽs�s��H�~i��
�?�%AKTX�Z��?36:�}���	�t�b�Ѥ��[Y�{�l�O�f��z�]���e�zܭ�SD?���1�쭇E�{F�5���a>�j�J�Y���g�B�����wO�K���w��&�p4%.\���|��:+{�7H���W��á�l�Ŷ7�b+\�+����V�}��_$Y)�t���QH�	��g�X�	4[�����[���h�<�ڄL�q�39�]��$z�Z L'ds�q�����1��ìC;��P�0�o�AY>BW�q�����p,Y�z]�w��"Oߡ�a�X+�����C����/	῁�Z�?�����w��L-O�J�l�_T�|���S��	�\��e& �����fh9���
��yl��J=�М\�V KW�H[�bk�Z�0��J^S�3�3�w�Z�W�s����|�3�Z"lq�#o6�M�N|~��E�r.d��[TF����yپ}���ޢ��x0�J�O�ܞճ7w��f,w��[~��v�q}�|mkO��9�������)1{v�_O��ɚ��뮵6.����R�u��|��/�2}�y=s����UV"���}�ߜ���N��o8�MV���^L�U�HYkl�_�-�&�O]���D�W�:ŭ����X��l��c�/�w��&����������/BO�,��iΜ�2��뼌�-�x�Fߓ1\�<�C��OE�A�X� �����*Ox	,��2��A�����g��c9Jȸ�7v`X\�]z�3+����g��h,� '"A��7�� �&�r�;��;d*�9��Ww��-�M�27�9��*��
K�}�lֶ�M�٣�׬T;FK��:�$�ش��;q��z@�Z&9�F�|1�K��	"�|���E��P%ȁJj���i���D��,�`��P��2Og�Y\V��R��&�G��I|��=Ҋue�8�#m��	2m�a���.8��V��k�qU�e4���9��4P���Ɗ�?�`[��h}��,� �P���-�
�Q��e�����d:e$��A�1�0�P��P}1��/L<p�YPOt�)i�<�d9����K]�B��&9����6�ܒ�i���%�Z���%��XJ�^��Z�cHR��uN�X�;��5���N�%.~� �U�깮*�#K <�N�x��e&P��;�*����w�f��3��� �1���*	e�a3�m�1���p�c��r���%�||��(O~)��9�Kk}tߛ(z�[T�]S�mH�"����TH� �Ǧ+,e�3�w�P�}n���S�&"�����Z<֛�ƛ3.4`��r�9�My����а���ę�*o6�T�]���4(�¶H�K�w��/[5xr���*���f�h�A�U���ޫ|Сe����Z��'�ޏ�
�N�z�r?�����v�'�/)W�^�xa��>�>�����f;��J�N6���n8�Kz�U���vL#ʟA?�nJ�E�Ɣ���O�N^�T{� B�g|��+p�t��w�:��r�CZ������E�jk5}W��/(E���ppۀd�F�����5��A��!� �U��jGo-�t��MBy�x��L��#,X'ڶ`�EX{�J㥮���IRЕ�`�f����jG��܏�L+!�@#��Â�v�d*��TWTf{�*ۨz,v�:K�Wf�7��jZ(zz}B�4s-J=γYl��_�Tw(� ��r<���0A*�Iрr�wN�;��-�w������L��1�����#���Muڙ��x{�!v���i4jqkPTqZ�)��!�{"|�f6w�/7#�P�DO|sf��Q�7QB׋�L�-~ZV������.���
�7$ƴ:#�,xb�φ��Ih%s�T�(��ӆ��賰aIp����$�a4�{k��EQ�.m������>�m�~�oq'ّ�0�\���2|�&Z\���̝�J����� ;#�a"��e�4��װOk���A"ix{�P^ŊGq.��B� �!1\vXN��ɉ�7��e�mSM]<�6��D��5��֏{�����B�.�\���l�lTk�H����7���aۆ#��;V��L��C������=K:��A����CsJ�r�K�L9EY��x!�zm�YDI~'��e	��
���|DiL�&P%8kٿ+!b��o�DyN|C����:5��}n
<U�x��_O9~�	�采;��A>�Ќ)$�i�s��>���dQ2�27�R���？��&�p��_p"S��*&�H���C�e������Ye2��`�����y<l�����h�{�=�h$��jT�e�?���۝ˉ
�~81I���_�$��o59�j�r8X��7NT�w4��Ӻ���Y%s?�#��)Tz��">_M,(\�I\Fۿ���|���s��m}����:���1~��hI���nmw�o��8�u��Q�c�vp�t�x�|�+_~ċ^Ѝz�ǥ��`<�K�s-���;%����vWٵj���t��8��2p	��j��Y�t{���[��8���זj�������F��J�$l��Sj���=�(��}�o�V�*3Ź��d^���q=�F=�Ӿ��6\�b�r����\axuF�ە��� y��V͎'�
Z#/r�A0� ��Yc�=i�J[xmrqT��g� ���YI��*�"ǘ�XĈ���x��zOp�\�/�璩�V�~�?𣻦�-K�&�M|3m�=��ơ��ښ@�#R��`nM.-$D����q�lUwj��u�WW�@(��74Ƒ�����Η�8wa�r8���oNU�E�Vۃ�e��M�{�s�gd/���$Uor(�Y��{n(�4)�ȋ����`����[şW^��v?���ű��V�0-���v�N2Z)'�n8rM��f��@����\ʄ��㺯�>
,?2��z��a�vb�P
�q>g/5��E@�G,0X3�v��f�)D��RNY��o�p����#����7H���?��;�y�ߒ���Y�y�\��ڧ��q�7Ǎ; �J��i��q$��߹�@��#ov�d��w��� ݕ����e�V1N�"z/t���҃$�C2�2c�#di��;Ie��f����(`���vO{Hl�����I�ë�2�s�z��Nb��nb��W/�mķ���7�����2pHg v���`�|s������M����QC�����-L��c/ h�浣�>NQN��,�xC-�CN&�v�%|���) �j�6<��m@8�N��k��jӨ.�e��@bk�=R��"v��y�ݛAxyG�&%Nd��4�	%B�f]}�5E-�H/�ӌ%	��U�l�9;=�`���-��L~Ba�/!i�b=(��\p1��I������xu��]S��/T�������
cu{����L�N׋?`��r1\�F��r
��8���ʦz%��ű�=w>cw���I�u�D�00�����\�Aj ��]��i)���̓��rc�R@�BWV`j�f�g�IX��X�9&"�x���N�����#_h��&�������wP�����Nj �C�R��������h�<��P�V�CAn�jBy��Z�u(��.H�(�Q2x����Ɇ�ə"K�P{�!���{�����EX���1Ə� {�pv���ч�T��sy8B ��MH���A)b&8�G��;DR<_�9qb��b��*Vp;�A��j|[g'`GV�1��v� f�D-x����alѱV��������כ���#w,�[���[������Up7�y�&��e��:ő���i6�b�Pcf��4�$�w����͒G~%pu�����?�+�E�X��!��d2��ཙ�"�=U�+s|�6�����8��[��$��j��IU�Ύœ���C�k+�6�}�/��/����K����Dj�f́"�9��ABR��d�Y;�-y�� #�)��S�{�_w�[F�״��zw��KN�����k
\�׉p?^&����_�%T�������`����6��P�q��>kr���R�\o%���P>���N��e"��ě��3_x�y����ra��Lv��N�5J �=�V��ZrU������k�"V��,-T1K��f�U� R��>��'��n8a��@L��m������T�}}���A���� �ʹG���Z����YJ\W��(���������������o����$�&�q)˝��5[�bs�e�h�Zx��=�֖�(�v�k�,R�%o�����П4�K:���*}D'��eX�2
zy�s�K���}%
K�#���*���x���i�ܐ�	�la�>7�[_����n!c���K!����y��Mb��iGN������ze�I}Aő&׫�v �t�������&��I]+r�1���ޖq�@T;y�+���������6ӵ�?������dF80�-j_䣮9/r���j�v0?�.ZQԥ�7�ɒL��am��#�[����B�$Vn��M �6����^~��A���$�>�"��Q�%���;Y�����k�>Cx���o�3@=����ϻpw�"����x�2��Iͧx�(2�I7�����}�ym�.��E��P�X���p��[h]��pA����<����2g��5"8
n��K��%�t��3f���S/cfd"���,SO��*;0;v=>����o W���n����p��$�Ϣ�a&G$�ln�>�hL��z0c��������aj�ʹ��k൑�`эLZ+�k_KDs�'�`�/%��U�
ǉ$�bO��f��9�d���#� �Q➠-��.q��!6gD@e��-�E�EE�ե���/�����T���_>YW�$�	ꢆo�o�є�����
�?o&W�*L�V?9�ه��5ޕ\��N�a�
��L�bs�ȣ����VX�w|���-=:�拏ۼ����Q.l!GB-�,?1����+��}��X�!��JvM�8~��%���;�5��l0�3yp��Y?�*��݆TOuǀ0�-��g���*�..}<�\ߴ�~Y�
�V�%9b�֞���0e;��q����jQ��n,�P�G4�/�֎Y�g~�3LWgo�
rlbp�T�Q%�W��e^��췥��d�eK�F�g����g�"�W~ЮG��\A��}������U�1Κ�Ѧ,0������qG��y?h3�ꍲMw[�y}�o��2����z�.��*��0+:i�zO��?7��~N��8�S���>�W�y�ܲ*f���N)A�ʓ�9�d��R�9�1Fs�qܓ@�,��F�9\��)�����`>j�A�8�5��$W���g������,���*R3$�����ƶM[��ƭ�/�T�C��D�8g�!?,�A�	�	?�7��U#/���&Χ����ia�~�������d�Xo>���c��<�O��"�0o*tB}"�Y{���M�(6�T��Km��H}�B�LQU!��)�l�ɍ�q� ";ddi�;�?�dY��)��8K���X�zY	��5���J��2�ˤ���S��[� �>Z��V�aI�b��YA?�HɁ���^Ġ� >7��*e/��t[�Z��V?�tª叢&�:nu4z��+����Q�f�W�s7Sw�ʁ8�Mc�L��g3��)v� q�#B����m��f�u��*|�u��F�oB|U�>C���m�{Vq����E�p�Cs_6��G,o�+1�	-�	fR˟�����C�:?��K��_$-�R��n_�	������tٷ�j�{�%|�I�2�����iO� �3��Н���O����؀l�xa�����h�R"O>ZiS�}����� �z�Y2R�6D^K)��[�E�X�FN�n���kfMm�`Z��²���+{OݵG�X=�ލ2�/��LNtB�廯�qV2��o�B5؊T��G�1y�6UVv.��K(��Z0j&�#�ٷ��Έj;����a B���)���N�K�hVeȬ�I��؞_���־��:Z�]����%QA:~�Afo?�&�L)��].h��ϳ�1�����\>8�EQYPT��`#��w�K�'���B��A�+%�g�����L0�(����4��� ��0�3��,�����GΌPO�#�d�.��n�ܛ�֏\�'s�Q���4F�V�����A��ҙo��	J�/�r�� ��jOH����	rO(%�V��fO[����:�U�%c������������˴���3]e��E 6�GO5���w��P�u��D�g*tiv@+���/IȌ��K��C RD28u�R�(��qf)�nG��/��8%�"0�P~�����W�	���"V	g��kV�E��=�$�^�q;$�-�����pJ�N�u�pc���g��ao+&��,�<5g�Xpb�4u���K4e�����H�}�\WX�ʉ����ِ0��������j|��(@�n�m`)]t�}X$���>�t8c)�q!%������,��i����xl`R�&Ҭ�����sBK(�e�Rw*�&�!iS�����|��-���8��S�Hg�$��>\�d�O�^�՛��A�p_��9J���n��3�e�u����Ke�ێ�q�^,�W�_�K����p��P�`nuY�$ �퐮%�K�(�ךz��d�;%�!�������]�A�K�3F䌐ft����������J���:wf/�&j�P��흭D�O��fw����@���6]^wD>7k�y%�$�
�z��=�AՕ��A3�׺���U_Bd�pd�ظ�����-��[Rg�36����8D8aI?Ow�-�#��c����H��tx\3��,��J�UX���5�.$�3xWk��d���]�F�:��rү�GLx�u��>E�ۖ� o:�����:AӜ�'v�G��0/P3m��2��V3˱;Se��;+`WCs��>qW��0`��n �Y؏}/~^�X�CeNiw�b��^紈����!
F�2[�e>'$�@݂	U�n��=t��H7��C6�E5���	�z��Ţ́L\;%+*���_��"��wg"���d?]�0�))h ��3D��������Q1���|ߦ��7�4����Q~�Ӣ��M��O�>�n�P�̆^.h��6mƙ-iL�2M�o5��SB���?�ip\�Q.:�T��^�H�/�w�.:���2&��_����aV�->]��o�����7��\.q� R����.A���3�`#�����ӴH��'2�IuT=Ǝ"S���ՠ�Ä��v��Hׇ;���J�AiKN�I�ϖT��|o����<�]z��f��
����}�\���uP��kE��(剼 q-�݁��S�j[HڽO�T����J�D!�57~R}�t��)yo%�f�\֏����2G��-a��_��ku�N�|��b�������5�"��(�'�l s�zbκ���TN%��k�5��qʔ�;[2����[F��s��ȽQ�3����N��I&	��� ��>����p����Y��%^�S�Oj�{��ӻ�F�!��o�/�t�ޅ�.����-z.<����q�YpBO,�\��ZB<�Z��;-�Q��1�����2�Н3���Z��.{���hn��z�.�I2�]�g{�=tR/�3���p�`�{�\�9~���7jlnԩǕ��E���e�A/ȑ%=�˰s�� x;	���;�2���JSmƴ���E�k��-�]d�۽�e	
3��j�H}�8��/��2>-�>�4��W�Z��ά�_�O��a�3�|pnn^Q��%!|��6).J�헳\�*����#��C��wL�l��P������2���:o�ձ�y���l��U����Ĥ\�'��@Z�/����XH$S�%��F��*I��x{�j��Ӭs��o� ���Hy2�F������?ك��Ӎ�r<	�+�%ao��=��S�M��J���ݛ�Ǝ�(� :�.X�GEl4AX_��En���(S��,�����2�̧�"I���cJ%���nzl�)NiN�|��իi����}w譝��ň��D�;�I��%�SO���{8�N��3ъ.�p���Tw�� �R��I�7��Ƨ9�i0r��?�	�B
��L��܃�j�P?<h�?f��@9�O	LY��G ��k& ��Rp�"���!����h}z%�Yΰ����#�����_��|���������|V
}���ks�]��_l��{~��B�O�17i�4ԅr�.�k.������.H�T(
�e{�ܑ�$�@��5w�lm�v�Ւ�8��	���s<�܃�3$�l������RS��݌�&ONF�ax��CO��Oju)�F��O޶!�{<��1N&�׫�ړ�s�-ɹ�̢w�r&�;��c�3:���`��-
���i?)�f�y�����Z1UX��	N|&�m?��<�릷�Yx��Q����AF� Ţ�@���N�����KP�v�:B�n;���.bo&Re�A�ۛ�{��ի 12��A.��};IQ��=i���գ{B�'��_^����������#�z |]Q9��|,s٪I�������i>���5�#�q,����%#�c]
�:���/���DRڷ7�FIw�Ht��	��/E/
d�ú���W��=0�����.��DqZ���M˟���_���f��np'RZ+�j=�LT�Z:�VN������!�]V���Y5���z�~d CUM�K�n|�وC##{���=�Ͼ�2C�r��N���@L'� �v�	�ٰ��K����u�z��Ҳ�쫂��XTqF]��lB����BOd���p����yE;Ny�9A���k�s�"c/N����
&��yA�@,YΙ ޲��FW�t�{8ĥ�7?������f߁�;1Q�Fhr�!R������,�B�b��`9���i,<kK�G����zm��׮�r�g8���'�y�`���������wB�S���Y:��Ȭ[�c͌D�)PR�y���E-1���a7�^R�!�C�}���ޗ���� ��6jy��P�o�����z�7��L>�%k�F�%j�r�_��e��:����,��E�a���[9���1jv�ר�şw��X��
����Ff�d�A���A6y��L��q��������>F��c���ž����ݡ��x�t�8.��� ��t#^���lzl�법�]Y�ߠ7`䶖��M<����V15kޑ!#�a�u��1�ї+nZ?>��A�l����/�E2J��$�%��?,{������#���0[J�Ёh�]��+��hR��=������\������f�ac<H���Ifi�QV�Ϝ�g��M��1@�ܩ��a�)�D��j�n�����3�uU�B�(->a+a�'��V�9U�YC�1ny�=H�0�2*i�h ��$�N�V�	^qnٛ�(�����7eT�j��A�V>����<>R���B�U
�h�`*TY�F�%j�c�}���������_�CZT�1�ژ�ጏ�� ч9�_��,0������
�P�7�Pa����ڀ*\&97!C�c(>ڰ��g(~3�_g�Ǖ\��Fj~�#X�Nj��V7��1'|kmu��ԖO�8՟+v"��ZW���Us ѽhװi��G�C�C�'dA�����U�w���z�����t�*t�p�L܎N���Ջ�$��	�����pky3��E��{>�
�xp{w�3Z<��JYzb��G��<p�ǔ6Ӯ�!Ǹ���E:Z�eLBm�,�1#^��T T5�˄���^tm�#I�ԉ�K��ԉ��mĐ3k��Xe��r����f�G�yy-t(�kP�X?%�b�ɿ��:�G�A%/8:��w���yǎ���$��<��(JE�N�n�$���`8N���m�V7�im����:��V���ͻ��;���ũ[	�t��q֜�-n���ѽ�9�	��R#}��V���� *A��r����ʣ@점��D����Ҳļ�Z#�=������a=d�X���{�#n���O�Y�o�|2�s�QYx��61���/+��I�\����"�6xb�3����N)���\\O߷ ��j^!ｳ
���������w%&�!��jw�fʳh�J�o=���Mˊ`��DG�]�>I�`��o&P���3�jM���&�� �_��*	��cQ.
IZQ�]�%��ԛ5�g��S��kځW�6W�o��'�A�j�I�B��?V�猂G.u�>�[&=� ��<QQ��6=�:f"@Ҝ�e!���:��2o�E�!�P`5���� �[o�l>?����(t��5�����ֵEAnl_�E뫅�K���lO&���cf5 �����z'&ll�\��EY�'P���mH�O{������G�ԒGT�,Ї6��%z�|�}�ϝ����J�
���g��!��M�.	*?a�ta����`q4z#�N�E���1,��=`ƺ{� ��7̏�'(I�uTv��4k����U�54�M��x�K�㘱�5H���%���b�l'�k^D�$z9�&��)j߶��[!��`Z�+�9gs�9�P�n���
v���3�z\u;�I�"fxN(�_<0����
F��o:	�٧���Ɉw�b���qN'�q:K����Up{ܪ}�˸���	0���A(��e-qY�X�*�X�����������X��>ߚ���^{���e�u�{�<y]�߾G�����$��D�Qʷ�k��̒P�[���d��ލ� a=l�x�ց��g6gw-G$<%;�x2�w����%���
�a���t�� tN'��<F�k$��i��o]������]����>�����3�V���,�U�����ǯʱ=�L���k�6WW:�d�)b�!!�!,��]�_0�:�����1�~���u��Yy��Kfd�|s���F�� �(�^T-b#���L%��n�Ļ*R{��6~u�8���<sf�R��-[����=����vcO��a����xG��G�X�>p��{n�T���x{t)$ט�l�'�y2DS0���VCY7�^c�d�r�_oJW�+}R���$����!�j����5�4,����z�!Ä��!���R�$0b��u���5	�%W��*�������Bo�Н>QkBxQ��LI]�r4X�d1��^D��wA&C��Tr��%�e5�t�S���0)�X�yAQB��7��~����m~^;ڞzb]�ȫ�����Byu�'�~��]g#��v��-���
�d_⢞w�-d�v���~8���J�WWy�؃h�HSH�B��o,z����g�.�`D�6��W�X_��j3芫��HXpE�������j>4SGN�#A��>E�LJ�çP����O7���A�E�/iH�\
��4ǝ�-VwJ4�8fe�(5I���swܲ*/���(ο+��.I;/�}f�AL'�>Î�vs{a�zǜ���5��@�أ�a�2���RiK$y1�3�	�#o���x�v��H]�jq�W8�Q�� ���BŇ�5�x��ꇳ��Iw�-�|Nd_�ʴ�!�=_�z�1�`ԃ��Y�ŝ�����ҾI��z@�P[�!�J�+C{o���~M|��u���b�Gʩ����?`���󜘾7�1�,� h�`�I��ښS���rSp�d���I"�Z�����tޣ�\��n�%��B���).�7	�[0lM@Lɣ�s���S�G�&��wU:�m��9-���S��� ��M%���Ć�����Z`��7l�L��s���1=qP�G��I��� �\�^ٴ����t����ٸ�\�6GK���E���7Ȟ<>�5�7v��wp�	=���c'�T�tL�n�}^�׺e��QFVk��9 ƤP'7aЏ��>*8��k�l�ߐ� �ʔR������1c49���:\e�<�Z]ۢ��.	o�r�R���HQ���+/�@����T��B�oحY5�R��|@c����|���
��P��Դ^�`�#�R�A����2Q�<4���T� �V-&0{���vd	=�\槷J��d�_�mC'��B����9k�5���?���O���@چ������L�2,����}��L����`����۳I¯��E��)��x	��t�;�!����y�Y 5�[HMϢ��ɶ�?��$iC�<F�����E.��!�=-�Y܊�����a�ԁ^#R��S)���xv�}���)jzYuKJ��o�7�~�$�P]�l�c��B6�y�tFR$��V� iQC:���9�����CP��>�AxՖ�W��7�~D���X��Hã=�O���� b���b
<��n��m���ܺĳS k��&`�4'�_A\��{
ո;�A&��s�M^썫�zҫL<9ف�k~jG=|�R`���SII����;�#r�t��"t� �����:̡�ap�}��Q�mR6`o-W.?8#�x��![7Md"�1�0��uvh�0 c^!݃�1)�B6XZ�;g�ve��(��w/>�)o�����q�X����Pk�Q(V�S.�Y���t���jr(�M����?I����af-��Q&���4܌=�*s�XSԙ���Z8�K��82�&��y����0%���R�|�c�"j4c��-�IK̉��8z(@��+�����j�>�:[�@�3�abBlʃ3���s���omvu�V!#IQYI�1�1V.�Ą���º�r)�۴�J	�R�G%���U!�A�D��q>�ĥa~ڗ�HU#���]B��'v�nGZ��`�R�T���=(Nv���Q�.��$�K2s?-�خzK2T�g_�|�{=���(EA(��������]q:���bϑ�fS�\NSBd�\I�ǉ9;�]��LtY��l8A��'��U����/�(�:���i�X_�-�n�$��*��*�O���)*D����f8��o[�a��R�R��[&��r���47b��hd��1�7����o�@�M��-�^�_)@���F%�*�/Qj�IuD��=��m�1C��(AJ� l�sEx�lc�����YX�7�1�VѥF��2i��Dɍɻ`��5%D\�Ch�hC��n "c�<�e\����7\���8�u&4U[7��6҅�2]򠕅��<f0��Pđy�{�$�TC������k�4��X�b%���b�_�3�ľD�_�ϵ�R��jH�ﰊ��8���8w�(=G�z���/�\x��M�ij�c����d��~=UW�)�O����ς�h��J��3��@�dKײ�j8��55���RW���Q�'
(� Z�[�A#�'�� C��V����	�=�ƣ�JR���D&�=�¥GH��h������"��g�ʆ�$┌��Գ]�uZT�H��fQ�_e~#:0�8��|�kݦ8��%]�ҍ�}WEBB��FQ�gǼPshC��c�7�y8�v6\�8����@�~���P�5�ۣb����,�{`L�>��8���>�hۋ���<��dƋ���;�6�� K����]����'�l�aHvk�?�cw��%r:C�G����R{��)w�(݇���^)W̙ى��EECǲY����g��Ӏ�й�V��[ͣw���I��Y���Γ�z@'��_��
.'35(g'�w��ph�6.��T}ӕ|��q�bm�|���vh���_�m�>x�s΍c|ů1�g��5�R�";*�;��ݢlTH��F	Y��U%��HF����:{
�:`@b�i}Q�����Ьᐦh�f���2�K���f��+Ƽ�w�:U� ��qKR+�bE!�s��)7����׮W!Vp�B]f�*��X4��+��ZmvY܌(�Y�hT��;J�����J��$ھ������{��/��=g�f�X��ĉ�^�x|�{�M�G�j�ɨ.�zZgd�t!~|$0w�W������m�Y�j:"Z|�AMl�G�^��Y�Z�y�*/mB���ϱ��šn�=\�i1Z�ů�K��y�?�ju�G�ޓ�J�5o�(��3���Ƚ��:}i�̧���
�n�*�|,'=i�!ñ��P��W�Q��ǊD�>5,��? �O�.	B�gX��'WOH��A�t:����JȮ_�����~�/�Z?�r����	�^�̎�J��F�<47q���р�����fbQ���Y���'x�����y�S
�h[���Т[�
�ꔂ;�>�e_�4�f����0"���ʯ�=�����Gց�����cl�$��b��+�VH����@�2<{*:��zy5��wn�:5�X��`x������$!�sd���#��@����|1��t!�'<�)&��E�b�C��RP�~��%�ZLĆH�bZd�>�{�Mm��cAuq�i��@����h�h��~�j٠�k��)�R��( H�������	�⥾�ֵ�[��?�a��4=��&�"^�8�Ed�9�d�.�ra��5F:�++q�-���Wa� ���K�^�b�c�8�%���X��
�<<����sZ��lCL�'�����?��2L%��B�8S�k�X�w3�Ÿ�;,�f��j�u,�;���yU9΅�����&��?��D����)�pJ��Z@S��6�+���1O�h&u��Q�\�?�����;��(uq�����gp�d>���'�vj�T�A����Q���oZ��*%N���19�	�[�2�N��Q��!2��4��!��%���a�6J�0��JpTwr���!n�h֜�E���z���x�U�S�}���Z�A��&3�P��W���4J=��L�C�5o�f�:�_��]�2�$ص4u'y[B��r�� �M���$ds���!��P�V�<�;o����	2��)sN��-C~8>n��8���[ R��M2�k�R@-P�;�����Gq<b��ȩ���O)2�U���6)g�6��v��Y�ɯX�}�5>���`�����+�t�{���� ���#���p��D�=m���� {;�K��G�i�D���Ƶ������d�I� nʏY_��
��鈺���"�YlJU":;�NK)�Qt�=����1��L���e�b�gT`�u��Ę&�Z��Qw��h�A��C%�d���̣8n�͓>��=5p��qm��zxe�l��a�$>pM�x���e	{T�a�O{BW�9����戇��(��(\Jx�Jv�UfAh��|U�ҳW:F��-�#����_'��zb�����Y�̙�gJ�f-�p���U��1����	yF'� l��CN�v�ٸm�q}�y{.��_u�9���`zC&\l�������Ge$(�dJ��8��R�t�}$��<O(;�9�8]H���Sӆ�n���6���kn��~���*:�Q0��Pd�r�v�c$�/T�V[��yDk�˟hљ�Dc|oӹ����8f�I�0�yGS�rmh�����Nžʶ5��?=ܳ<є(�,�D��������i��NK�oяL�8���!*"f����4��x\��`�~���� ����h������I]l�`�����w���TZ����s�pԉ�?�9��].�@K��,�V�Y
B���J}�)��.���_!���rіy}8}�uxp���.yv�I��)=�4x�$����F�X�J�~��+���7a�c��^f�e����!S�|��R�f  �L�L���2�0�ܶ*ɟ�3s����#�`���Z�+ڧ�b�m�[�� ���&����v���5��i��@\��95w���m&���L�[�� tN�߇
)UV0�B��VD�9g�/۾����BDq��"�o*��z�p<U/�TsM�ӃM��jЗ4�yL�r�\A�TX�/��ʮ�`�|92�^��6)��[�y>�̞6	=�~�1�(��Mz6[�6�Ǳ��ĕ�̡�k�-��}! ڔ��>d�]���W-h���v��Z�:~n��!���U'�%D9�f��Z]�爮n՟E;�kK�js���B���[�0�E۲�m�X�o�ep�(��O񓅫��8<���&m=�]YS�Sw��4���2ޯl�E�b]Y_R5�5PJH��e��I��'��A��#+\�dx�g4�)&�m� ����-rN$���c���*[���aF�M5O��L���hF* �!�+�?J��s�M{n���Q���� ]�jl��r��FQ�&�G�!/s�7�i�4�*ؠ�[�򩍂POF���	�RW��صb%�Hь��=�éiݣ�飨����.}�!��2��Ϝ�H��ɉ���
���M#S  ���]l�f\ɟ<�ׇm'ڑt�Q=#"��:֎�Fq�� )t�L�8�ʪp�ᡀ=�Zc�5������0���鬁��"�P���%Z�1�aI;��y�y�����"P�����Y��M�;����2��qgt!j�M�X+�}���=J�͐c��2�T%ůg���c�$�rO�X����OC�������Ñ�%usa`�ᬵ������r����Z���]=K��&�5�KB03U8t,�~`����f�Q��q|�5/^ߔ��trH̢�а�C�-���a̅��ӹ���3j.C�'8��ɘ��7�_$DSI�5X�JDP �i��7-c���'�s�9��\�+�������z�N�=��Ux`����w&��|)��Db�`��;�E�Ey'��R�erPe-�R��Vk�$�K��L'��3���V#�M�RtnZnx���1.8�]��8��&+�Ȃ�q1DJ����|Y�r��A���Q�uW6�)ٌtΘ���gK�`m��+}ɲ�����]�s�L��Sbg��K%�<�%���O�3l�ӎև~dAH�f�|U�%�Q�'�˻���4X�ş	|��A���o�#0*u��!�"��S��*֑,��]�~�f/��^J��yX��pÒx�i��R0�
������_���{���D�����g2�E�5fHhH<h6Onk�)�/ohG���D"����U��aG�R�d5*����'���x�ܰ^阤�j%�Ш�@��{�i�F��݅]�~�i��R����%�4z�ڸL�ȝ&��~F��kC2t����3ۛ	�)����g��n�Z���V2˯C�V�G�5��9��'���0��@����o9���py���x�dw�I��Q�Q�KW�Nw�iW*Z@PↅP�yk�8�|	�L���(o��^Q�	��VQ��u�ka�t���F�6Ct-�>��(*��qS����w�����e�(��Z�A����c %%���s�1�~@u!v��^��5d�`)H�V��o�<�>�N[W�ʍ�㕨�_QS���Jdr=`fr9SB�Q� �����a8(X�ݺ�Y��п끗���L���� ��;B����N���j��T�IqJE����h�huK��'�Tй$#����~wM^��ǻ��A�D1��LJ�g�Qf���.��&�����ơ��V��6Z#P����L1��n��T���v	}�N���3�g��gʞI��ps�[�86Y�$8��֚p�n�2��V1�4[n�BY6/��-r_��p�����t+���Ӂ�Y��g��3�@y狝��-�[5�yV# ��A���f��T�R㹲O�=RQ��!���ƀb�k%�\�����cR�KO������4�o����'C$�}�z)��R�u��U���y?OI�Ѽ*�(Qy4$�h0��Ľ���L����VR�;=�9"Rʳ�����}��_�T��A�P{��kܜ�2=�ǭI� �i��Lpp�]?a �<=�
�;���Ϲl�[vr�"Y�T:�i�Ȅ���a��Da��#��:��\���A#jcA������UЀ��(���@1J*��O^���־�~�����;�9��vքE�>��]w����Y�uI��)sF�;�ֈgkj0P�L&�<�u7�:���
Np �P�D3m�ŝ�z@a�x�	د��/�'���̮���d(s��R5&2&X� ��6#�Ik���y�K�S�i��*����$U�����
�?8�%��#I)2�ӣ{f^�{��B���ĺ�>���`S�!;�3�{_�����꺪<��B����1fQ�/x.��HW@��^�r�;ى�@:�a͐��`�!���c�CS��a;��c� �_�e�/�afi1���F�8ԩ�Q�Z_�0K�}#���
��I@�c����S�u����[��E.�Uu�44�_yb��r9@�skd���҃��["�a��%n��^��.���ܗ�������4_��΄t���q������5~���A��n��K�F��,�rw��cPQ��VPFF��+�V�z���jٯl%�ͧ1�&&�2m�.5�1MfvJ��}��&~�:9*�?0[���m��xI�ZK��S@��]�Oc&��!
H�]�����͐Y� *�����I��x>�^IZ����b�e�:=��.�[��,օ+��Y:�e�m�����SS��+-A�!��0Ǭ�N<��;���\��B����x��SQR�;�MFDL��m����%��rfnuR �	�Z��=l�Fz��[<<��jUnZ��Jd~f֥3���oKw��YD�R|2b�B�
�������ݐPǓ013yA ��rvԃ.�n��o5P+��Xg ��)�ϝ�m�'�Dl�#��P��l45��:��Q�B e���q��jǪ��x�,�c˓�����q��OB����S�7��-X��Gx��Չ���D*c��('ǽҖ
��ʹ�h���h���{���'�͡�C���l��S��|�5L}O�؅1	��n� Pi����䩂/�H�'	Q�����{�N"y�hS�:�s�%�{M��@9q������S�%Z��h��>���+��#h�cE[�5O39NNx�����ƭBb��{nP@���_f����C�yQ��9 [��4��jb��|�:�+#�d��("����1B�!�^��p���;B,\1��IC�O�w�Y�M���������]�� +��а���n�HtZ4n�[c	h����t3��w7�K�/ޭ��6#+�(���E6��;w����_V4,.�b�����4�FIŷ]��k��,��@�Fs�?�|��,Wؘ({-��;}�\��3,o�<�ro�A�n��(�w�a��\3�k���?���qM�k���}i7"�'ڰ5�A=57��~t_H��&ȉ@Ʒ�J�۩�Yk�i�h�&XK�~^�[�
r�DE8r�Ln���3����ƌ������$	>#,����&�P���4/��C	�'�t�zr6��^S}J�=�M�K���]�c��O1�Ӈۥft>��l�2��\������̦��iC�����o��#�*�K�rk�;��1/{�اD_}�`7�GS�#�?~i�A�7��;���s��@�E����V'�N>g��Ʃ�*>��� ��To��C��!�qҒ|����M�A��ǋ뿊�/F�7L�on��"�$KD�h7K���E��v,���)a%�|�3e/��0c8��
�'����q�h�Rp��	_@�%�	��K��ڤA+G-x%A߯Ά�^�tw-�R1��H��/5�\/!$�� ��"~J0�qh�{T��uft�=T��b�����}��|��B��	G��MUK�@��a�?�nA�:I��z���8�|e�CP�֢��o칐���>^]��X�n�I�Ϋ�	�wGH7%��y�$�AU���˧���rֆyCP �[���Yc�'�G$��ba�d�����n��?n���D�6��`���I��g3ig��G����b���=� ,(�Վc��B�J+�Xe�&���p��vV��x����_*34U���v`v��4�(8�~���:=�υ��v<,�33-�T����2���w�0�PMNE�zՆ� �@q��'�P��/���1�朘�⦈:)�oOX��������Wa��1�>�S�٧�	����$ʭ9�r�/�v�p����7��&��\خ��HR�o�7��-�ոV�mg�r����X�� ��&�Qj�:�������.z�����23g���}�z�4���&�̱���=}NL�d�CA�R9|w��S�Z���_>��:ՃX+���κ.? �Xd��>�L�y�ۍ�ɜ�x���^g�<+���4u�����0DGNm�(���-V*XA�+�߫^d�u��#���W)FL�=H�ݏ�*$	��$l���3{�gf����B��쮵�s'��Fd���Yg,/<�f]0Z��^|;������Yq����\8Ã���^Ƣѷ�AF00�5:�{��E wt���zJ~.M˿�њ�9��h�s�T{�y����;`O�x������u�4��l˪\/���5��4�tn]4�:�D�u)��3UZ���s�Wn�}h��d��x���������ob����Aʬ�������--�M�~�<����jr�)�.+cR���}���rG&�pGh�C��^.����&'n��2(R������Fۺ!�O���p�i�/�$d `���T���N�f���^0��d�m�Rkm�O���Y)�\��P��{l#�0m���0Q>�>�LE��l�b旘U�c�ۍ0�$=���O�u@�/\Tt hW��u3�jZ�R�E�5�_:,�'�Gv
#hYZy/�`���Ů���_�1e�Dd�4i-���/ɡ�0�)��u %���H`�7�BB�%��4��Ca>`�uqKp ��I��}��j�![����3<��3����Ф����6���A�О�U���?�}���`�c��@���cͶ]׍�zo �8QC|��ނ�h�c�ʼW�p�"I��2[�$��05O�Q#�{T�%��wd�D+K�����-�Jg
a))T�`H}��]U*rlI欷�J�Z�0��Ջ�YZ�C��
HG����1���ȍF�UX��$��=7��+m�xa
M�[)y������xh���ʹ��c���2+���f�WP�˧�WQB��
l�H@ep�U6
0�]��ռCRB
�(6���!���,vLN�_�K���8����b��^���A��y�Р��y~N<��`S�̟a�����)X"V�:S`c�������k�G��u�vR�b�9_��{0����5*7�U0#��!��K�"rs>_�����Qg�ir�-���U��w���(�5kC�����kRq�y��19_˶�=u�<�JZ��8:Д �
�Ge�Oz,���(���:cֳ������	bd0�/�������LB�イDZ'�L�R��)��+����.Q�E
�@�6�S�a�x��z�����H�rh�ƶ2(:�=d*�m�i�ٞ^rj%��B���I(C�[��¬5�3	��{Yx+�G���;�hp:����@��a�.��-���j��9���-9�{�#F�'A[�;�Ś�}�9�988�]�*��K���x
�����G�$"q/��o���jO[��R�F�P��n�j�˵½�����'�j�����Zt4�nBM؝�Mt�{Gs_9�nN�=�89�%x�V^#k!��hX��_�g$yl�X�v�P?iC�6��S�.�n�X�@�^��u0��r\k���V���sdp�{A��Lp7���rn����r�U�f���_��	�-1QY����+�8N2_����o#,"�_<S0_ը����t88O����j`�C���U���=_K���TUVBg�շY�y�����=�:��,S�6�'��Z��S
��Rr�
7�+���Qq.�:��G�y�.�A!�b���EYUP�}�W��h�͈Hr(�͑��`�����kya@������5�2 � ����/��ʤ�sF��C��߀��� a�1���EJ�z��w��iL��;,�9;ƃj���z��b��FOcRBg���n����?��b���	Qd�aVu�(�������C3e��x.�M�.�l�4Qi���uƩw���{T��Q�Y���"k?��VJf E�6�u�'�挎݁Z�'+�7��v�<w�������e����G�A�� y0�r�.�a���!�x�MR;ği҃��[E˪�c�J#���D�YZ�`�W:�V��f�~�_+��Bz1.�!� �x�S�r�uڴ"��2;��:\�i\��'|�s�M�[��Q1�ei�n��q�4�H�<s�E}�1�s��n�3Q��Y�t@�׽ �io�v�`x;��a�5Y{n�����-ؔ>��5DSl]��w�4f��foٰ[0�v[y�$؏X5S��Y�8]�N�a�Jj�[gu�H���(�)y��uM�y%�#`�s�6��	ʨ-�����Jn�X�qKg��vM�q��p��mh���rԳ'�	�5�����M<�]/����p�Ʋ�\���%��=}(1�b���4-����2in�t�QVݻ1����� Gk�/�s������^���NBo��ӿ>(�n��3[)�� Q�,C�6/|���/%m�]���H7�2ҕ�LĜ//�-{������lDw��ng,��f��ּt��k0�W�eq���=sU�?0.���c����qm��ү�QC��S��᧸ǂJ��#E�.��uz)��7!�K��{*�ŏd�k��wP�c9k�ym�	a�;oAE�L#��/nöc�Ar�C�xf�^���b>"��]Kw��v���9� ?b�@��JfO�V<���2�d���l���Y�
H���_N����E�&��f���J[�0o͈��H��xFꂡe��6��������"�D�H��U��H�����|�O�=�EC������O�Ȳ$OX7d��ìnl~��B��|��yG�p��)��?����/��d`����/�<aDx��Q(�iN��U���C;�<Z/M�೤�R�L� >V�KV����7���Hd�U����w�d+\��_���.ݹlV��!ʾ�"$�8$@sS*d,)���c��۫�^�0\Z��#�;^��F��쁆�U�f�i��u�.�8��{ .���2�x���8s�A�&?�B2i��C��h���h�k�d�P.>����3m'3�S�F����Ĩ�3��֦�����C�ָ��J�^<�e��D��R� 仍ݳQOy@R�����9�aN�����@�I���;J����	���BA!B�l.��#+�-&|9 ��KCY���9�"�x��b���p�*�+� �z����{��+k�|,��B��ײ:�F����Y�	0�#+#�~D�9U^�J�֝��.G�-� �E�GIa6�a/��~���Ӡu��F{��.pۉ��orE�ڋ�?D,Ј��d�G�~/���X�y�Z�O��.?w��R}�����N��ep����aTօ��n3�XO!��^��<�=�[��w^��/*�5����V��DF�q#?�hh@m����n)9`��d>��O$]���%SE�Q��1����2l�#�fsA��{a��_��N�w��:,ؠR6�sK�f��~�7ڽu��g0��%�/^GF5���{ A����xf~�D\����s�����b$f�uyJ�̣�,B�z%Bt�颭6߳��7\�G�B�'�-�0���Wg��ؘY?eBv�:x9%������������E��	Wk�?)`��v,'+O�Ǝ]��2�d����c�!|H� ��YM��؁Qa�#��f�0�������cPa���E��,�� ��%�*nkI��|r@��p*Zy�~gN�N����6�y��jzG�,�E��K����ںcׅ����x�.�/�~.5�Y^�."�r��v�<q"�����l�p?N� V�5���u�@�p ���|	��g�.N���he�T�1�޹Qc�sh���rSޫ�'o�w��F;��%��\�.��(]�G��r���ۧ1u<��HU*-r��o0d��6�I��&�K3��B�lZNA:�rߏH���!䬀�ц�g_�G�fߔ,F<d�8�?�s*�ؼ+��M�W�ԒeBi^L��|������dM.�	�I��k	�r��9jg����nPU�Α�k���7��׶9p(7�T�^{�Q�q��i��e�.�4�/� =��)7H�z̥�e�q��[���ǘǬy� �\0/�I�X�hg����Bǯb.����j��e}�@p�`o�R�i�������%�,��)H/�=�� �ep�H_TSL�,����؀���cgP׮n�Y
�D:W=78=�`��;���335�}��Uf���i��q�
},,mՠ�����;DO�k���w���=]�}7�v�p��a?L�N��!�Q�l�l�Z~XO�!ά�
t��W�f|c�̈�Ϋ���+�K�O�:U	�"�~���#����W�uo
��B1�����1�H��u�Y�r��3�,d0@^vC���1�iV��h��D��n��vd�3��h4���%��7��ڋ��n)�z����Ӵ}L��X�Y)R6Y �*	���}�:M)�l��$7�#��~�՛�6�%��vX�F]�p�W�83L0���2��H�왔��*�^��	�4O`+4���)���y���gH0J��q���mȞ=��y�g�*�����B3�c���^)2��bLIN:�&�r�dE���P4�o�KB��A���\{o"��M���̓p��]��$��4\���0.�0;���qor>��!�3����fƧI���B�7If��x���<��U�eA^�jA�� 5�J�}2�9�9T�;��5������n*e>b�dv�ŧ�x�j�E�eE
MD�����4�7X[�[�c2���G�q��4t���dz���0�]Z� N�@94�զ�^^����
2�����=m�x�P{����j1W,ӽh�8��.�R��/�\��d�ٕ�>��`9�(f���t��n�(��/��כ�6��Ђ��G<���E;
��6��S�����H��	�	���E�f ��5��x[��9v(�S��1G�3%P2G3����dV*uI��؉��Uj��I��ڛ3]%(�Y��1E"�g�8C���_�0��C�uZ>h�8�4�\C����ز8��c��Z3��py{�H���Э�/��ߏ�Ǫ!q�6|B	�T�Gk�:��;έ�q]�"�?�׸l�u��T�RWx<C���z�knf�mۧ�na�����%^������:��|,���A�jZ�dX�	6aYb���c֝J �Su�i0F�#;��0��z���We o� A$Yߑ��J�E8�Y�F|�F���0�������޶-�M��9�;ͽO��	���-�ns�#1���ҭ�d�����B��>ޏ�#ȡft�����m}�X��ٸ0�N��ay���N�B-.�<�>g����~f���r,Xy��P�v=�eBo�&y��Bx�.z���׬���5��-ӣ^?u�6lqqd�O�^X=u�Ӊ��"�N�y�9٘�Q���\��
��a�C�g@�p��,��<�kF���86+��L@��r��GT�k}�s�$�����N�w�A�U�J-��DV�����%l��?G�����I%�%n�Vz�ZKF��U�,�w߁Q�b�?���)�^��!1�0�����3ڠ@�s�YS�q���K}���=����Pw����X _Lw��Ǌ�葥���' Md�`��24C<@�
��8|S����ŵ�	z,h���V�M��L�
��,�JT-&�n�~�A��*��j
�6i-�F�&l�
�; *R������KƦ������
8?��ٲ�-���Z��Pw�75�R�Ҹc��z ��]hK�L�lɑ��g �d�B�r:��ߍx�W�jK)%
%Ӵ�����m�h�����3{�ˊ����M�e`q���b�`6�xi���JGi~lD�#�0�c|3몍'�X���&�t���o�z�9�R�@����O�l��(S�±����9=��������e��
�sB�G��$�c1�9퉕��q}��m�:��*Ch�փ�Dͅ�ǂ?eB[���gW�~��˛.E�(�׸���o�D������2�� ��<�	o���R�a����ꪆl"�|���a��@���W��Ri{ԅn��a'�&`�w.��W��-���\T��?��ϥ��Fr�͇z9�����("�3��"o��øۺ�@�O\�p���^:��K�dޒ�f�#�2��.y:B�Η�:�Dz�U��T�2t+��\�-�X���6�
Bw	��QE����U8�gѬ�.=޺� خlݰ5>��0|~b
L[�j�+eM�q�+賫�����+����=LN�NbO��g�������s�"��tѤ3(�;6H�Bt��@��Ú;�H~;&�1ꔹ�Ƌ�'�b�U�Y�_E:=�8wm��ųF��>8�F���?\�@��>Xwؐ��~���Vl��)��D� $��b��4q�tN�1��X�,��&1�Z闹u�#}�l�ɼ��G�2L��X���/��!lןSLaǳ�8h(�娗Ӈ$�e�#a#E����A����a�Y��c���c� ����f/5Zd������猒3��͍�ct���4DV1?�R�x�$~>�2�,wF�����#��PF*�I�-+�8=��_��%9� �;h9gqd[�2K2�����@�gO��>d;�:��vQS7HvYy�q�!i�Z����_��]ܬG �ҿL˿�aHG����(��w}����	?�ܙ��.�=ﳧ1�gFx��N���b��t_5�D�b+��t{ʻlQ����sv��������s�&u�ɍ"�����������?�Su�Rs��A�u�au���i,/������E0�:��Y�	7j1��m�/B��<��%xy8RGKg�Z\����]�k�ݪ��DC���Z 
� s��x�%iB�y�h��b����|���L{L����%&OKr>����1F\�2uS;xP�[d���q1��x�}c�d��'�:!�r�� %�pf��c��N;R2C7�hdEya5����m�b9-mL>Gܲ�|H��o��K�T
�)B��'��Bv$��U�q��b"{��.y�RF4,�֭P!�ڮK��B���Ok3f�n�_�+-d��!K@�t�2)G�sd�JtZ����ֻ9��=y�|ɧ�2���������+H�:�PФ����L�ݧ�Ja�����Y[��N�Ȱ��/��SZ2�a�o�f�Ӄ\�&�x��������G�#w��U��Mx��*��?i��.<�J�O���Qm�ؿ����X���<���d���؝ I��U�{�@U�h��(�55z`ƚ���3����ĉl���}k�5�X�o/g3	a���C�SS���:=N̬Y�	q�<�
J4Nf����}I~͖mf�
���������8��&�GO��SE/"/�u��F#Og�A}	4������1���계6�t��]܄U���`�f�ERK1�?��
�v��.�`��M1}�ტZH���#�4Je�#�S�3����¾��o�����nod��ަ
�CY�Ry�h��s%�cR3���gz.7�k��[ ��U�k�4�Ê��	����f�<�f���	���?�݅{���]���r�l?wc���OP ���5_���5tp������^ l��AfTF0I��>���Q+ch`���T�ʋiA�d�i�������J0�<���oyԗ
�)WB�ړ� yy}/N���y/ĉđ�E��'���a���E�#���q/�:b5d�M�_F�\D&�@��Q��WV<Dr��u۱��C�[�3�)�w"�oDߕ;���O�Ԏ*��Y{�)j��f"Ɍ�v~�����_15��LU����n)�;�@7.����2m���%T��`e�j��Fm�ݬ�B����&Ev�EW��M�	M8�y�#�ÉH��V����?�.��?��-Mw�������5J撹Ӝ="{�Ǣ�NE��'jR�\�B^v����d�OQq�#|Þ����>�tNN���uh����瞨�0�E�ؖ`I=}�7k�"QU�ͮ�i��pj��l��{k�c�f�]a*
�շ���p����KJQ��L����s���@KT��:�����E�&�!���ZSpQ���#�愥�����ܾ�`�O3I6[>��_	��m\������^!{��O�aA��F�V���쳥#b;;݆F%�1��fOɓ����-c?�)mo^� ��be-���x_)��}�W�Bz�2j\�rd�ap;Mt�a�{ya^�v���f/��P�3FF(k_���8v�(���!� ;7��[��#�l��������D�>�� ��� (��O�\�zC�<�󻃦^F}m�jgt :�'�V$̘]yr��FZ��^sL`�P
w(��m����U7̓ȸ�Gp�Ʃ�5p���6� ���M慌���ceD�^=���g�h�L��^l���&FlR�Z��t����LF�.%:�KD��GӄƉ�[E�{x���m��t�}�^>vu��ua:ǩC2�S3r~.\ ��3`�O�#����_A�v��.�Շ*��Bq���ɒ;?9LL	�m�*���3L�����b�
j������@(b��^Ӑ�P{�]j�p�O�h�B��T�m���+��X���ɼ�x*���ws,^���p�RR垌=4g����+5����@*C���s��_*%�\@*���c+�l/i���ey{���(`���/���ĚRsK��w�F���4'ͭ���&�	�N�(�m�2Ft/A'r{
��}��@5l� ��=>4Q%7?!��3,�+�^҃m"�hh$�4���pP��jdWr�[H���薐����	�}�����$4�݁��`����w��?u+���p��|�c���Y	�5��;��69JvPW�9�|�J0<Ab�Ѓ���M�Q����ϗ�C��/`u�P�
�	̝lğ{��'X? jDCQ��j&�V�_9���Ih��E��,��^~li!��~LD��6wlkj�-3H��OKf��/��nB��w��E��25�Z��9�O,��P�� f��������B����p���:/�t�@ ��"p:H#c�7',���7<�2+���m�,@4s��H]������x��`�a���?���Ԏ;O�S�
�I+���+��Z�Y;N��Y��h�����+��bEȪ��s(��W�iq�=���5�mA��G�7�ݾ�Uf!Z<`&�G������ϙΓ�?�aĿ�?f�s�����	�z���Zt��5�Ҥ����I�hOs�	ܰUT�y�i�|:O�u� Y���m��"���p`����[������$^t�֣h��w�Z�����N��%�H�Wv�]�ł��Ty1��ܤ���H)�������ウ�uv�*\�L���Y{FE�C0�
B�����R��i�'"ۈ��n���.�G�h�G�+��3IPn|��#@���[8�:|)C�G6Tp6|��۸v�/����$E�y6��)ȹ�ހ�?��������rV���U�l��5����׏��ǋ#�����B-����ҽ�5'��-Ft|AȾ��b������t�[���F73���R�%��Cf
��d���	�l��H�l��uTJ`T`����4H�q�驤�wG��x�dI���*����Å"�)���H�3����V�ˮ�s�����zR�/�U� 9AQ��-�ʒ"^8#�a3h6���\��}�N�`����Ji��C���M\/�k���G�t�W��︠#��@�w`:~�w�����$���ڐ��Ș��/�"o����K�Eh��c@����X�����@�f^{�h�Í6-zW��Ǹ�=��N�␑R�[k1	����Y<ҟ���8�Za��8��R�6l(�n����w�K֠���|�wt�cz%�&��\	<�7�p��T��8������(��"ͅ��0/�Q�VВ�R�l�"=�*o]j�d4�)UW����!��_�~����a��<����[+�v95�(혮��/��~Vk
9���O�;�]��J�nVB���d��l�m+�j�W����.�a��j�m�鼶��au�I��	�(�f72�������;hzm�a��`�!*�k#5�����+�3?l�O�B��߈Vz�p������Z3_u�Q��s}rN��SN�ڛ�-��cD��ֻAR??\L1�	ѥ�NǸA^	n�U����$���w8����3����KqQ�ϭ�RnGh���[=��A&�2��И:-CHц�:E��~�3���]W�Id='m��v#r��!	ݚf��Q��u�μ;�Q#cd��F�~��s^���]Xj�	��K+y$�L
���R���ϗ
�ū���pN^��*u� h��B�:3��p�e
�ۺ/�c�wo��̈U.��0hݤot�������M��Go	S�r��d~�d�|�����5�O�O�{��9��N�>��Ilg�w�y4���3��TK�-�W{�H�|h �Y]��bR5[b����Y���m�.@�Iӛ)���=���c-��?���e<}/I�\��Ҁ�|�+�ZU���;�]ó��ܢ�G�Q�j����ij%����bR���V�g㗡�\8
�5�b�P�������҅���E&��2��,���A�DJA6���	����ƣ& T�3߭R-�9��<��XYǵ\Y�ǒThIR����d�w�d�j�R���e?wX-,�2�#�����k�w�-����t{(����»�m����<�K䊕~X���Z�}N���o�+O���%����DQ�%�b
��C��]���%a8$��{9�Rgi���m��!a��´||8�d����P��f ����ׯ8�XC[b�kb�u�Ol�tИ�CP���G	qC7�EN��{�p�[����'�NY������=?���c"���m�/���j5��8;��W���1o�nj��c����g�J�9����ۺf�ա}SY�>�>�t-����)�-|�s�V��,�1����=�pV`?��1
�$�Q�X��*0J���ꐱZ?�~��:��o}]�i���A�=�oGt��6*B�>N��ʵX�"�2
�w�g{K*W�K��cvj�
	��qa0��:JE&�o$��L4Z1�����%8.4���1���=q(��k�})�j�[�T��C�,��Sq��� ;3���z-������<y��R��#�9X�Y�O���o��  [
N>�Q�D^�&�$(�m֨5�Y�\8/<�gMөny���v �2�1�Qx'�y{��\�#����)j@���mnE��[��)&u������/E��� o�;�Uj����C�E�
��[0
0d��v���$�t�mP���V�������z����q��7�^t�0�@4�QX�z�0n��M�j�K]���TL0��|�}�a�JļJ��T@5�:�|�F�Z�$�CY|ŉ��^��G��k̝�0��!�WP�,
1�r��։7��a:Q�/)���+�e7·�/���v��
���lp���}�&{u��U����PkP#�e��w�4{������:�hr��w0�G=\SN�/�������=���*q
�lh3J}j��c�*O05�x�?avl-��{�-
SS[�%򇾒�шG���`(OJ� ����5,�5o�>���1x�;D�*d��w������(��٢���ƌ�8�Л���IRO�:��9AG�n���$�6]����#?�٢�z�M�T����ݝ+�~U�E*��si��uf1
	F�JAY�ڤV�u�}M��*��04z޵�:��{t$�_�9>�� �2IG�q�^��� ��I��v�㊕g�=@;D���}�Rx�����}�Nq1�Y0 H��%YO�t�1�$�
��$~K�ݦ�{��Xp�2H�4>2�(DU��MC!��1�,ڈ4G��\XN�9Q���E߼����#Q@��E��(�x�u����58̠��v�y�5LS��|Hǚ���x9V��c&Z��d�n$��lE5�N�w����f\��m�1�(��ixIY�Q��^=6���0E!S�:�S�W�<�� ���n9傠���Z�MZ����J�@H,2���tӼ�>���eHi���i@��J�e L��e�EHO������Ð0eb��3fChX�z�|o<��O΄�#'܊�܀qb�:���L�|B����%�g��O.UK��_�N�&9U?�C�I�3^�����;{r���+Q��N?M�ne��Q �����a����0�t�Ӌy�AO~(�X�kk��i��3	x��9�W`���˨��p��� *�Z|y&,�Ij�� �u����� �����0��Ɓ�J��Y��p�DKZ��/��}\C��XU���|��p����%��'V�۹����+�K�o୮�`�K����!�أ�=|��S�Y2��sLQ�z.��.^�I����Ԥ.Hz7��{~������2���C����`(���i���5/��[|��N b�}�.F:{�9�5���8��;.��;��I���CY�L�ߧqV��^ڝ�6��٦�󸹂Kj��0��i>�L�2��!4�[ F�Ӽ^"�j�8���'_�5�uN���>���eP�츍����~7K Am;@bA*6��Z|�n���j/ׯ��}�Wkd�e��G��H�K�׸�*~@#�k�52K�u,?���=L����薸�
������tQ])^4]blj�*-�<�����J���'}*5���݁�6�5�F���c�tnŔ�𥘮XK���6��o
��<����0�M��X��8g�K{DR�4��@Fz�/�r�&��rB�э���ϜB�����W�xP�œq�s�i�|���D]��/���>�w
�):�Ɦz�J��ڥ)�-�6#��o��hv���l��/������m�C+���0h|��8�\,<>������[��
7�Is��� -�o���உ�w2n��^"]Ꝑ��- ����1����8T�W�I�˗Y��₠��:�D�_�l�mb��~��4$�'�ֺߡ�\���9]4��E��O�u燨�;^�#�5FN���X2i���'�#��1!ȋ����ժY!�:��2�=T	9������[X�m�s-��
M=5Ԍ	��r�:���L��A?5��>���Y��'bܖN��(O���y�`�z\?�{X����a����h�h�bW?�����@��J�Ȉ�u������6�:i������m���W>�obH�1�=Ls!�Y��I��t�|��^��l=�;$в3�1�2�A�G��t��n�X�w�������Ӻ�S�#���&����~�,m4���u��"I��s�I�u�}���qmU%�>����S��S��lT-�J�V�<{A/��-M��p�����u���=���sx�s��@��O�4h a�j;J�q?D"3�q��3eYs@|�	du�y�\}GШ���UPG���7�PỞ��;�%��4g�C��:�`*t�9���'8�m��u����q�mZ��e�T���j�6�p8�f�ȦY� ��r~��)!U��	�c���\>�����'��\{v�����(G<G����3iQ�����v�k)(�rn潆~O�� �=������/oE o���<�(Y(�s�*�<�\ܤa�@�an
�9���U�mù��'����̽���R���n��[�ʬ��"VHÜT�On �����W��w�����j����&�!��W-gv�Zn<��T�-�D�;�񙡂��OZ��*�n�&0��������(�m���W��c4�i��k�#��X&f��Y��+10&�sNdlq�yoZ9�:�i�.����R�6��Ə'+G��Y8����mQ��@/~���?։o�*D�~��3|���NQ�u��<�P������d�}
��/�������"P�r]V�U���m"@N����4$�?*�� d��kQ��K/y�j-�}o
VV�ώ��� ��ʙq����EH������:G��>�Dr<������2Ou������,�׍���ɒZ�^�^}s�-Z�kjRS��pJ
���W�V�);�B�� ��r�%�%h��e���Y�'�=)��u"릨��e�V�k;}���&����=�A����B�_�0]�R{Rp�԰	pe����5!�%xC���5wJ�"���-bUM�9�p]W禆�b����a9� ��zެ��Wog��7����6�{Vu쓄����5B�x�`b�ɮ���e���6�XQ�,n1�m$�r%���2�e�\H/�����y�eI`e�g�?�D4���@\!R�pX0��T���m����0���^�Z�b�sq؜�{�Xby2��xaȴ�ĸ�i���]�YW��V{�W�J�/�]O����t�ϓ\������v�����A�&_��TQ��xg��f�C�P��N�*������	������I�ܒ�&���Lp��R��.����r���+Zd�;ԫ|ʷ��7HW 2S�Y�c�?��6�lXք%� c5����u:Q������7m�=�J3
(�t� ,�u��h�eBֺ-Ӟ�4u��ٸ�{��x�m��*�t�-�I�u�I^�s�,+ekMl�%�:��|"gW��V;R���d�3>�o"����+l4�����.3���L�|>94�[":�~՟�f
�_��U�e|��.>���4�,��O�����������|~W�����:��^J��Fx[ �K�l�ӈ�D䚆�tzM����k�6ug&�@<�i�:BJ[^��#H*I�����>��@_�.� 5��f�1I�����/*����P����t��d�W�O��a��-e��F���.I�W�[I��G7
�a��ܩl;��SQA2����G�~xH̩ϥׄC.�����H���2��/�����RN�TiF�Ă뼜PeK����[�%7��7�z��h|�I�c��K	0g�&U
��No�]�g_e���E���S�A�1�еT,<hd3O����E����e�w��#?��g���hL���u���z��ʕ (	��ϟU�����~VR�qZc;��\И<7�#��q�^a�����w�)Z��X=e�:�&�pUr��}���C�D�C����s����Ȗ2�֘a�"+2z�v3��<@��h�����Gg��d�Ͱ��R Iޗ�ҷ;�6�ol��G,�?�s����9��i?�y�jH�Q�;���ր���Hj�[y �z�C�}y�j�i�LUZ$����<��H���k��. ������۰���_�r��^���#"⡧�$��k#�o�p�]C�-?A2�}��1�F*I��>��ۿ���*�g��1߫c���s��_��|̵����1�F�T����񾃌{�%���g���3'È�� �%��ߞ�%P�kX�E�j����/ߚ�x���JI[�ӫ���Y2��*ǾW#��g�W@-i���fݔ��\˭<��Ͱ��<]��}���� �i�ޮ�1��-�f�|y�W�Y7y�ax��ꎛ�Zc��O���e�	�!l'���븈r�o�5]��ڜ�I���	 +��}J�XI��n�YPd��4U�3Om��y-������xfu�zd�����d��c5n��/�K�#=@��=��߰	��kdo��fD1GW�q���$5���4Y�ϙ�oo"a�9�ߺk����~�Š[�8f����dt��u��A��C��e�X�P�9?=O�I���l�hd���0��h�?.?�I/�$X�q2�A�[�3��r�Ю��>�"@�P��i����[DSo�
 �J�:���I_�q�A��6�kE/���r�l�R��N��dS/O��e�]�yn���x1������;���;pZ�w���r�+_3�ކ��Cز�q�̤e�>��">��c�rX�m@&�:H-���oǸ�1x�yr�[��g�LV -aﱢ5���k6���o�t� n\&4�ٮ�m�-���.�1���	�^��7b5SϮ��m�� Y,�������9�x����3��J��\�{�K؁�������c_��"�� ���;��Kފ�-J=.X��~7��':�xN;|����u�'Ij�Tk-���>��b�/Ǭ4ُr����	8���u�)��av���s>hy�EC<��S��2��W37\�#(�}�A�߫�� �4��MR�:A����Ԏ�¼0��o�W[ s���M���\���w��z0�����zut��J!n���4J��g`P�8�x�L^���)��hn/y�jI�Ik�ن��aҗ�H>��o��v�r0_�|�5Z~[��	~�v����X�hM��v0��*�����kVOY<n���c��dL����h�K���Ū�:jeo�;
5%�>*B�{{v�Sb�Dc���-�{�� �]v+�J��7l`�X?�M��b4\���]��w]�I_��Dw�(y7#�, �Y��x�z���ٹR✚^�Y���&�:�����e��ۅ��G�nB����^g��E��Y����6����Q�XB�s�p���%��<�V	b�
(��C��� 	E��M�	�ĕ��o���`�U����kTV�T�[@��˶y��H
��	H�\Qܛ�&A�շ�'�ykʠ���M����
＝� L?������1�`�Jͺ-��D���?�2mWbn�[ޜ�v��Dz��]/N�I�I_�ĕ�z�w����G3k�ϥb���`�LW��NK���(@ׯ�4���W�B�y��8�n"U�Bg�ﱟ��yD�a�� �?�YL�ziw3Z,'����RWL�p���g9��/Y5����]/
��V�>� ��e!^@d�D� ���L��SQa��˲�1�#����2��l�Lk�/�i��b�[�I;����\�M�e�g����31vpц[|^�{���}{���ʳص���4�%����K����M˹��WW��6?�TL��PpXRyi��q	s��o���Z;�#9�4A�Zz6x>g6D�DCm�������Ϯr�^n�������R:\F��.��9�^��/̈�ʉ�yw|Մ�?�A��)9�34�ؿbh4T`S�:���u�e�WXc��C����siJdE�N�����6$�6��QA-��ω '��H����4���]�E���R�y����hF7���+���������殳�t�>�5�$Ӱ�D�0Hf��^!����%�ꂋ��[�D<B��S����/����8d�;Kf����� 58�����ޥ����"n�E��Er\]3���p�?WS>,�C0����nиc�����E�,�zq}cnn�P,�*��
y?◻���t��z�0���0�p�Γw<��>��qB����4(.K#,�]�6�EV��wN �";�c ���x����Q(X!A��o���B�=SX������O3��Z_��J�U�+q:���lb!�wv��s��RP纞F���%K�s��OxEoz;4&��A�O¬SO�?�~f�s���0C�L���x�θ�HJ1��$�k��e���>Y��x���S�.~����(���`����iۡ��̭d�C��

[���v�d::1RS���ޟ�O�ۦ��+��u�:.F��4�=��/ʝo!�l��p���
��O�<�ƫ2��Ӵ�f|�j�0�8q?�L;��,���s�
����O�����y<g��z�8@($D�X��s��*X��Q�X��ّ���\r�� �����Ԏ1S�Q^�-������{o�EC�F��h����d�!��Z�����뢦$M�R��:������PX!9���e�_��z��Y��4��:���a{y�hr�E=}��)+���Prj�k-�����=(3��v�a����v�(h�P�L�J��?�)fL�U>	�g��s�s��Z�B�/�_��!�-�ԁ��Ov-�w��JP�JĴ#7��c���X&�ܸ�#UM
��݈�ɑ1Q9i��ZB��ֵ�a ��xP�3��b��~?*5�(����6J�u,�<�e��<�cb��Fd)?2�")TV����J�ҭ�=7���)>W3�����e���j��>��)p���t��(��ҰG��Ks�{�\��Xq( >3���Ӽ��Q�5�d@W�X���m`5���s�5@�
"��+=ζN�Bz�U��!�i��s+a{i��֚8A��}����5��?DXS3�'i�E�`�T��(�H/�SD��Ɍ�c.1�ۗ\�o��r�̢��D`��&�4��.��G3��u��Q�A?���]9�f�����WL�ŴۄV���Q����7ȵ8Z/;@�T�U̒��1���}液V0���4��i�_�d�q��˅cx�K��~�x ���\�\���1T7@߈�W������l��D�6���RE{�Rd��Y`��� ����u�Jǟ0��+�m�p�϶ҏ���o*��"��,��'��:�M_u�
׳%�s�1{�B-]g��N�ipqX��p�0�N��uQS��(�k�Љ��*9�j��epg_��
.�0��w?Դk�t��?�>c������� ��}�ۺ�C �,�5˛���Rt��A,�,ߚ���6�/�Gz�0�<�T��H�$3�����2��پ��q����,�zq���֑tB�O6��1����T'3�XZ�������t�s�_�0�Ƒ;��F�U�@�Sj�=qdܐ��e#n������yYn���*�*h5��C���b�4�ȓ��c�s��=y���cyYGq�`�,�J�=	͙Ů�zH߽��� �b���k�����Y��×Ie�=�Y�WV�[�*��\'I��Z0K>��`��YUKn��Nk�=c(^�g�>tlɝ�~X4�d���?��Mg���YZ8!ֿ�-�������O�
6 �%���h� ʙH�������+���۲�)<�z��q޾��x����qW�Tx!�p��UҪ{���g���huP��*���FB��]�
�~�{��Fm�P�iP���ҋ_�3�E�-��H�����-r6�e��`�E���!#�nS�;��Us�a�����\����"�by��s:�7ҥ(�v==(t#���Yj��Ky3NS���r�m˗����ՑG=!����x3)4B!jٯ'�R���FRfԁ�8�A�b���4����1{K{7�?^��q��2�I�;VQ#��5�d����ٌ"��d����s�hw<�rx�h��L�U��x�jg^�_���,��\�ٯ�����GΔ��|~�%9��M��0��k&3f
4d aa�4/ ���/�_z	a�H;�M�~&�c��?64s��f�\ת,H��X�e�IMDߣ�&�M��_6�S� dp����fX����,�����y���j�V���T筅X<�-xJ��Rݦ���L�ڙԽw�2�z_E;Y(_0���TT�*X��k�l�U�Ԋ���`�!Q;�];@Qb��+!�8b�H�"��x��[\OG���_���M�yQ����h#,&v����	\U�d]�����Y�Ӂ�1@�X�$����z���k����.SG�jF�.�Ab$�`�N$ȴdُ��X��	?ql���wp��*�f�H\������Ӄ�9�R��0u[���a.HM>�	P�㖐��]���^��8^>�ۂAgQE]�$�S8�������=��&hh5��W����S���>����XSi�NFu�	�<`=2��8.nT~��>E��mGXMv#b��H��ͧY���J��[|Bܣ&b�d�_v�t�p�1_��Љk��O�sp���~��M�|u�˥q�����mM�~�@��s࿐��է!/��O���[m;!	K�S`�L�ۻ	q���s�#��-�֪t�f�� 3Q�m���W8��Dm�A���݁���S420Y��`S�-4D��w�J*@oX�
J�~r1&7�z�prI������ZʫW[��"(D�E�n����?��Z��gr�m1Ö3=sѳɘ��"�D���Z�H��xلp_��M���=@H/��%s�'qB�ԑ�CwW������h�ql�f=�K�	�&�_/Yb\��q{eb��j%:�_1�x�h��\��AA*�\���_2�ܞq�Pٷ�VQIk�l��� ��w�)&��v���`����c�t�]"��g����z!~O���y��S"-r�3��ï�lNv�0 Lu?=g���Q���u����^b�3������X'���|�n,�ZPk���[�?���e0A3�G5V8y��m��)lP�G���Ia�3{�$8�5�����t���40M��M�6ږ�N���'n�k)%$u�kb�y
 ����D%d�p,'}���w�*��"��a<M?ap��(�L}�LAŋ���!�d]�u{HRw�T[�H��xOL®�k�o�����'�x���A{�m�����r����?������x�$?�������PP3m7���J����y=:�P���2�V复�Iitc�$M���]�Y�Ƴ�P˗�̖��hXƠ���d�l�%�@)�.V��� ��dp�>����wV�rߏ
�3P^��⣤�cu���ւ���0^L��6wj��.˱���l)�fT��ݹ1�W��1��7�7�3��|-^� &��	���a����Q���P7�Л���ȉ�#��N~;�j9*��<G�i��ZldI��_�����O.��;�B�S��"7�8���n/�C��Y�aM%|����~K�|m=uG���U9�.q]�瘜�)7%��=�U<i;帬��V\?�m�c7P����C%�;�j��:�D��n�A����$�kd��$2n,������U?�� ��^�ՑU
�q�������ؘ��h�z~0����9��_%���'g��[�7�3Ѕ���4Ԩ&�)���J�r�;Ĕ�R�K��TѮ�/Ώ�Xh�7������$�6N@�#�O� ��0����P�fc['Oi9H��Kku6I�� QM���i�W3�h|��l�q�KlƆYDh�R����t'P^��]��m�/x;�z��� ���T��ۙ�"�;����<��¹��[1 [�0���ƚKl�[*�r�u�ѻ�Z�3�iײ.iWO��=�Zh��d�YД�.M��l�y[�ƪ��rG��G|�$����euF7#l��14m2�\ѪJ�s��O�=0�O��:qt�F�tG2�������-���*�ӵ	IAe˘
�Q�@�'q�"Nx��ڮQ9�I�w���Q��N+�6�����/�+��b'(�W��􎅕�l)������u,�P��:�R�T�~�jI�J�	���%ې=��x���(G�?r����x�������p�?N�T�X��R�Q]{��V:/�,�{N��c���=�����=AMP7�����#�b4BIl!�<~��% ~����߅Sڑ��y�ݗ���N�x��&G�a�\��h�Ƹ���0���Qk��J��;�������3�:/��� �e3.�i�_�ϻ�R�WxÔ��c������3B=��(���	FUj�QPל�a���j�F�Ab����[U���&�ͧ�f���i�� 4��a_#n�2���Ӎֳ�H��a{���u��ٓ��[�(�2��c�"��_z��9Lf4+� q#�5"9�+�^�,dm���s�DiH�ꆈ)�p��Q�y�η���ta5bL8���]��(��«���a9� ���&A1};{�U��.�
����:;���Ew�"���g�Ơ��?R�@W��@��T�x��[Q���Ή�}�D����SA-s[2}�}��>P,�nX�.��1��q�v�ͥM��}����֙F�4[�a��z��S���Мջ��Ծ̅����ǉt�42���Kڝ�u�G�[$*�,�T[�i�������m�&x���ip*��I<3�'�8ԋ���U��	��b�������P8��H��SJI�o���Zb;õ�a���Ya�L����v�7|!hf}h+�x?�q���_ms%$�h��ּ��&Ѷ��caN�	C�l�y~�v����(���4�Ib���e��
9�:�F���`9$���I%pP6�<Ħ�`�5s�i�f�y�D��n���]H�ζ����Z���1�j�R�bc"���w.�ZY}>�� ��>�$*ć����؝��j&�6�'���9vN��4��%�8�r���w�㕎�W7{�@�P`�	��6�p`m�0�0#0s/乁}u�9��Gx�'}���ry'3�[0?���P���c�S���K4�T���'x:-�R�&�=����O�jO�{���]�3诨@u�꟤�Aݥ�4�6�b��/�Y�k�M�)�FO��}qq
~���u��Q���yEI����p�gXvU'ox�m��)yq���.�i������k�ࢣ-���˗�y��M��'�p��~�)��-���M��6�?���8A�t���B?�AL�H��h�F[o�N�䊚�7H������s���� te"ޢ2&�Yqˌ� =\7�]RrSd��:.�A���9DC�*Y���9�Xt,Q��� A�Ʋ��:�_�+�
X�T�
'���?�R�Zs�_nG�R������P��Z�_�~\z�������`���J�3�&*��$����Ě��ǿZ��RoYBF�P�
̠*\���x�N%!����WS �,�1�3�ӫ�^��M�xN�6�1���������_D�F�`��*g<�J�tc����w�LڶX�ۚ�37�\�B#�wUn��p�aZm��_� r��l$�D���[�&b����&7�c�]�yJ{s�������͛��M>��tj��X�.NٰZ�H'`(���1�#�n0����������#�8D[�.�MP3��5�X��Q m���d�7��Ie�Q�4Ņ��L��8# Z:����LpZ��9��@��]!���4�xa�p�j��#�N��������Ͳ�s�U8�o���0���]��*�Y+��L��� PT �]��-��2��~��r�ɥ�;�n�^g�8�ag7�
�/呮���'N��=r�����y$�e�%��'�)��V��CT��.%�����q �_���i��-�mP�n���.&����[x���FNڶ_Qc��S��@յ�#�,t�x�]@rr�[Y7�z�q�B�v�L�X��Q�X=��E�(~�l�+��aZ�������!,ucUV���w3�fベ%��h4�ߒ�?�&�Rb'����	�Y�ʤ�����ʢ����`"@�I�M��GMЦ����e���" �ݏz��J#]��G̃�8�����C���~B���?�H��7qd�$���}���m�U=_%U��K,�h�Q�8�S�0~y�-&f/!�p�ܺ�zՅ&�=�d?~��T-A�F"�5ـ�$λfmޠ]l�#v�����]�ŕ)��������$�Z%T]:��<Â��Ԓ���(�3!y	?;eZ�8i���"���&Tv����\����������T-5i��������`��ԝHL��bD��}?ȥ!|2md]�f��K���x���	=�C�M@`�L��"���5����!Z(,ĸZ>��Q�����b� �oT���g����A{u�ڟ�a�*������~�jy�e�����m��V���ىw0apPo=���ΞR|vd�eӪC�����"��9����FWs)��b�;STx��G��˾���E�l�j)g��DV���<��~�E��}�������Ha�� ��况�o(�EA��G��kr��4��3˦�\��e%Fe>"���̭��f9�����@�S&��mS�x�M�*t�57z=/���6_W�V
X�57��N^�����|7{TpEK����N��R�d�h���WمͲ搿'D{Id&�@�,��T�&�1n�V��݅����B����ĀCs���iW����4��
�լ*A�I2��V9迒%q<�˓��v�.V�E�;�:B���Q?C���R��f���߭��@���l�fѵc���F���1Qi��	�6Z��Y3< ��6{6���&��v�N^��ٶ�Yjs��%�2�p���Q�~��@� ���
�RMK���)��F��������{�56����KG���ϲ�;4X�l��G�J�je�B���I0���֣5�����ⴾ|c2��������F�|V���r�_��;b���0��Bu@��b4+a�����L���,�?ɬ�!�Tx�~:�U���=�]������6,I>�&��k����󈣣�1�ZM�+1"��Յ|t��t\���I��>�y�y��	�a���=Rã|�̝/���P�v*0����s`C��:r��4�<�=zk"�2ŋ�RN�Xg�"���G:- !���v��.�4#��MR}�y�7�S@�>8<r���ȶoI1��	�r��:�`fB�h(樌���X!�D:x�ߡe[0RɮQv�y�Dp/��H�U�}��0ݱtģΥ@������D�1�_z<s���|�+g�4��2A$� y�R���T��Z��h��\P��MoJ*Qt��\H�q��3=XS�m����Hp^/G��A 7Uh�sB ���pf���;��u�_��Lp�<����Y�vV��iL�㡬Qh�:1L���_D<ԭӺD�4��C��Οv�K>���l�IY���	(����~�G�5�1 ��J�3N%�%��R�3R��@c��nL=4�-r�v��΅����ۨ�}ˌ��#0���.�H��2�%4��N��O�x�S�e���f������ Z�@VA!c;�$1�pWlw�Фd/�'�ŢD��kg�އ>c�tz�^�p��N3Z���EO�� �_z_|�<������c����)"A�`�06��$#�>]�%ö��/�v��#�"(1��њլ@��&`�"�z�2_�������-��#�!���[7q��}c�L�2�^��5�L5�Lأ����B��#�ѭ��)X��ѡ�{�1��<��3�z�=���xZ�}>��`�y����g󒃶3��P�E�!�R�A�q��5˲��y{��\L���+�����Z\|T��`>I�f����5�I� �}���
C^�>�X���Nn���ee��pgA�$��U����##a���!M�O����4�g4���N�~�δ�v�k����o�w[i;W�}�SrO�/�0)�ׇ�Ǚ�p���S��uRG���2O�Bb�d
S�����ҙw1��,�(��B��������`�.����J
@,P�1��E���}Mq�#�1�*v�4K��+�v�����`�����B%������[��{*����}\�	E�ͬH(<S��ɺh��Y�e�.Ž�[�E�b���!s���w�ǔ{u>�vPt����CGE$�@DL�:�Kr<�r.;�=h�z��m�d�I�bR���.0�&rI���f��*ow6�V��!�\�����Z,��1[ɑFJ���X3�H$�k�.�u�/��a�ob����03�T���Uo����PG�7�qg)����\d�u_Rx!E:D���sM$����Q�1>w-�e�K߉�Iؙ7p��}�%yi��ӝ1%]�������u�?�	��0ͤn+��ԃ�ϱ�����u5�+B��\��8���>�˓��� �p�xl/�S�����*�>��Ĭ�⨔�"�� �s�@	�]ɡ��9-�m�5>t����v�'�!|�6��4�eʀnT�]3r��<ǧK��ώ� 4@#;��U,R7��ʟg$wF�n~,j�et
��I�=#���/���� 1K]���Čj(N%��C1��{=���E{|�k#V���.��*���v\x%���Լt��t����?�|#�EO0y���0;�O�VL���c~��<:O���^1�<խ�z�o�5d>P� B恟�����X�~��A��Rg�Y� B��(ۦ�t���Q���-��w�P�/_��J����I��ƴ�fm�w����C�F�3@8�=��6���^�|��í��<�>r���1ZFM�|�k:o�=�r�7
�����Q�	D���4�|�7���[ T��Ӯ2L h�R����áX�@Kd6�(���D-_�!y�G���"�I�i���	����G�K�37��mS�u�
�7!+��p5������sIK��^3z�k�$�|���B����B��n��Yc£�Tap�c`v}FV��F��%��/���j����ZN�#�r'��&Pm���g�hyS�ѝǨU����?D��sۑD����jɂT�������u.����Q�=�J�*g�հK��C0Ll�Gp��Z�Z�$6dS��0$��U\V����� ��m�U��mQ��,�"��m�j0�A�C��4Л���~������5H��R�U?(�������10
�p%��O�/�:�1;Q�%�)ܥ�¾��%��@-)U���.+��D;]Ӱ&��LyY��jM��hҰ.NYs4�0Ä�b�a$�E�O�����m����k�eY��d�0I*M˹���!����m��&���law=�s��*����cվs����!{и�6Zh�d�X��˪E��{���Z�M�) �=@ &fG�)V7����`TS������������?7���xk_�%�a>4�`ؽ�\�J��57�o��/��k�![�P$�y�+<����W�� ��q����h�3>�O��P�N���~����g2;���o��u"gh!֬��x���3���όşz�"ɻ��N�j�Q]*n�4��xq�n�K������tK2wT)F�2�4b�ユG-jo��W��7@�Qv\��W�<1pUu�ǴoO�f�9cPQ���7�uH�P���W�u@���ʾh:�Q6���>b2G���۱�B�_���ީ��ƪKҿ�n"j+�cж�ך�@}�/��فl
2��^ѹ����_J6K�&S��ϛ��y-F�-���JI&8�b�^(�K�V,������s~T�DoWd;�̝��V���L6��|]��8.�'<&��8dx� ��uS]/W��6��J.")3W�*�L> �R��hF�8A0`�(x�GA�{:z?;0�ZM�+��/Y�����З'�b�S�"e���]���^����	��|'�i���K�B���I����f|����cD6�T�T"��Q�F�a󟃅]�_��&�{2�w�7�y-|c�F��~�����֢>��L��imn�N~�[B�)C�x=7�`^|������̞8饆a���K����hq�QX�أwF^r�%�Rj!����-`Z�i�7A9Z���B�Af�?�Us�c�.��z��WE��8Tњ��R�}�����N�X�*�A{�#�ޜ$T�*���^�+T������B����UAE��·�����=O�5�U��z�����0w�m���� ���5Q��@�0k��m���(RC\�6(0%���1�}�1[�`h�2��n�LBՃ��Z���T���hհx 45ëiǣ�)��B��[�Е$�A����aF�g-�8,ie���1���e����X�	C�R_��0�[{�/���k`=¤�TF3�&�g�Y`�	��T1~��3���8~�Ӿ�.��t�v���BL�����L�ȝ�s1�ʴ�9Cр^G��(����1pynh�D���p��\T��+���9i���Tj9��30-�g*��5��h����l���q�/����	�<H���:A3ϓD�BO`��(3&M��6"F7aF�����})��J��D�tk����2P�9Y�Zy|�
�w�Q#��A@f��C�[��s�<�Ug�?�7Ш�[�c���%u)���-�s����7��-"j8�6	��.�ڨ�X��������rF����=�j��U ��#���1W�'��o�MT�H!�1�x��w�MY�(Ce�Ȩ�q�u��c��ѷIm:8%rm����c���U׼�v����,�{�e���y0Y4������'�X�2AD��J�shM_�)b�����6���|q ���e�K.g#��$�-��pG��g�����p����vo���< �KKixâz�I��� U7�����xj���D����$�2�^I�`�!�.g�]�:]��R���cD�S����\���rG�b�L>�{^$��(�B*=���w���/0���Ě�Qc4�2q�P���]<��gڏ\ń�(A����n���+��)��^P]w����u�ZeY��  ���A���*��t�{tm�O�/,���2��#��6�j��b���-9�2�Mt���򀴱1��UR�@cBو�ù>��ey�D�L?�P�䩼��#K8��B�J��ٳ=]>@r����H���O[O̥� ��F�Dr ���<'��@ڇ�v¼�v[܆����� `��wV�1]x2;(�NaÊ"����B��އ B�N����̎����]�N {��hr��1OR�8�7	ӽ`Ҙ�LK�ӮRJ��Q�29`�6U�9�Ni�S�>Rݬ�IKˢ�M��5�$ˎ�P�B	�_Pks��Ms�^`o�G��2%0+���kZ�|aݜI�)/85��u	��_Fwq�j|o_����N�%C�,�-�h��41�KWA�����C�n��3�M�aP�� ν�^�f�m����7�*���Ryw�L�=X��-FK�{�#�4�0�-^�3�m�P�DF�Twȕ�s�bc��Z)�����bs+�A߰���f�_����,G�f���<�����?|!J���ڋm����C넞��p. ]1��ra�'��^E���g��$�
'��m��E��am�g����K9���UŮ�!iV
#ȠF��o]'T徿G��O��p����w>cuO�wbc!����BE�i�tA\��x�W�66�R����Cp��qa�r9�i��)za��E��u]�5{a`��Ds�ٝz��>z&�8��!�K�'���� ?_4q��AQJW�u����i��?9�}�eW{A¹Ë����)O��^l5L:���!FU$$���� k�r�%Y�Q��.�wC~�b�@}Nm�ψ�՟meO#��!��^n�D�����D^�ƫ=쌧�
f��5�@�:����2���"X��R�~��u�FK����v���&�|l��h�A�6����P����Q�{�GBa|,������Z3�z����mo]z��Ɂ�ط��%�ä��sTNF��P�ǘQ"���
�b�����=�'�����AZpՀFy�U!S��A���H��l+
�xc�5>�sG5�o��i�pS)����	���2I���|u��U6t���ү��"QŦ����ׄg�;Ju�|��v�^|tW)N��I�EMm��uP<�Z���c�܄��xe�r�[v�+"�S#�_�ma?��|I{V��b��X��E�;Z�0�)i�M��s���:+�ۮg3F�8����mD�oU5S�lm�0�6d���C��\SH?���Lѳ(��V���Z�� ]� KCtp� ���k���mhC �?�oC�!შ)\�.�+�$�(�8+T�`�X��w��u��|�����rd���'�"�M �v�yL�5N�΂�]�g���;�\�3!.�)�d�_����� )!V��Q�"��Wr�/:P�B`�h����O^y�F��r}���({���:f�c%���&h�{��5��8>�j�%~
��n��l]4l��}�NO���w݇�ЊJ�fVl�n�c�C�[Qᘔ������eR��X���R,�r-�h�;`�A4�B�f�>���TBu%c1z��� �wE�F.�E� ZH_:��m�� �;G���|���2R/όAߌ��2;	��H;�*c����x^��[��ڦ�(���@��%>����S�!��0f�0#(<��#��bh������j��A2COJ��j��* j�3l��֋x�7s4��M�tC��o����Z_%:�>KX�ā���|��b�NBρ�p'�,T}Tv�N<�~s�AH�`�5��t[C����I[A�(G��҈�g�ŕ�,r����JCh�>A���»G��]��	O�,���ae��m�Q>�-�ت$�L嗌�iH�Yŝ측��#s#��0v�?s�e� ��.�F����Ol3�T��"���<+G�It�p≐����}�����������}���m�����Ŕ+�0��Ԙǐ�}rt�my����-���)�^�X?�Ù�ٟ�� c���!�A���9���i��4�{!�]�3>�DOE��I�?��Q-^K)��m��5��~�h�	�hA/pP��^�����J��O��+�wKH�0�=w.���qU���F���<~6v�#'�,80�F�G�?�����R�x�o�U솃܊6�KJ�����a*W&�����hN</\�{U"'�6Ǘ��L/1��M�H��ڠgB�Z����Ц
r�+q��h.���E��)�r��&�c���ћ,K���F&��:��oc�ۗ'��U6wT����z�Z�bB�U��]%0�z�P�>���S�@��j	n{ѦY�` �U�< o���erM�s��jq�����i�A����t�$)吪p� S5�3֗�j�S1���H[>�'Ӯ7u�ݛ�r+m�}����=b�����Yw@
��;��:��-��R�N�st�I�S�%�<K�2jܿ,�����ߺj�a�k<_��z����=�V;�j���q"r<����e�L��K2ѯxz�殧�s��	�֧Og�nr��#ޤH���S-ע��K�o%� O;pB��c+N��d�Mٲ	N�i�+�G�<��E�b?�uv�ϡ �H���5i��Sֹ���5n<�4��]�G=�F�N;y(~��p�I��qv�u
���/������pK��T~�*5c�Q�R�d0)�Ɉ1�\@w)�w�*��{�l�Gp������IҺ��əɤ���=E�Z�>}�g�c�i�%/ /2$�rн�x���4��g�Њ���`e/6z?:?���ou�v�u/��ç4�x����N���� ��Р	R�fFU#��1�MS�`�0���ٱ-�Z�+��j�"j�N	���e��M�75���2H����?��C�Ϲ���1��\��� %Ҵ�΢ⓚ �*����F���L���o�lh����5^GWLf�[��=�rňf�`Y�N����3@�_@�-����J�"�i��Ȱ��cz9��C����ژ�%��W~���1{��W@�載/�C�ٔ��x���33��<g��zT���ɒg,��PҭW��ς�UHϗ�c��_C��������{��q�nT8K3���~�-��j+��ٶ�v�����dtsH��{%��9�1O��;<�[�7�]��!�f�z�4-n�be�i��-f�FY��+���7�h�i�}5/AKLG�%�����n�s�𘔱��'�gR�¢<i9���If�I��<��g$v!��M�[���-l���Cy��W<���Y5��������65���P���KKU���˅���q��K~oE��e���F��sC�&���짵���Z����8z0�(�Q ���EQh>!��h��$E�����,����\�;��Kު�@���1}�֙]x��9�� �NY��#X",�QN֕��_�x�zӶ��*����=@M�"�-ڴ��{�?̀$��_Ǡ�[�����#�;�ͽ�J� p2�[��g5�8X�s��NFe�a����g �c�6��ʝRK�W|��;�U�M�c6��x�MYY�%s@5?�vnC�C\���Qƿ�A���7��pY�f��Gڋ�d����š5�^{C?�Dw�K��f ���j�� ���w�(-�Y�Z���ay�t��5�+�H�*�q��qyQ�ϕ�V����18��3xS�)M�}����@]��S���,Y���q\�V��t�R�h��۱&�Qi�4?<����_��~E��KH��'#�����fw��C�J�iU6E�Q"7oi��[l���xo�G�8=����USy5B5j�颢l��	k6���r�,mg�_��U�͚@zS7���D��Ȝ�}5Q[Z���P�S����4SV*�
csPa��G����ۻ"0���\�F�$H���57�#��;�sC�V�s>��=�{=�X�a4]L�0�->�D���a��Fz��4�ǂtRa�%�@��SIf����Z�Q*{�<�7�)�1�N��Š~��7����Me��)C��r��&$�K�viK�2�&-�]X(^l�O�IZ�F]�R��އ����~�"6���:��;��w�c<�9Ky{*�; u�]�2&S!��-R��t��	R� C(�ym�)��:B����T`�7�wPZ�)���E��[�����_E����xq9'0�Z�=������n*oo�1����_��q?t&Ej	j5Cr���r�ߢ�BRiF��M�;�����Ue���)��k|��p\%�$ ϥƊ�Me��׭���r��]h��N��\ښ�m��)���z�P��Yo���7l���.�0��gW/Y���>�^�����Z��}�UU���Q� Oto���Dź,��ψ�"��$J�%�SY��>�,o������śB�8�����3���~:��[�xL��@[ԖS��V�s灣���=�~� �
�U��p�V��-eR�0�p���5����+�^2|}=5Le�H�tjX �v�Q�rA	�|�.8�?ri@֫Q~(cS���}8�-)X���33��%Q:�r�p��ŷ��%�]�"�tm����pFĞ%�Sf�	�
.ٲ�Y"+��&>-���sD�I�7rs�e���[fȺ�s_��X�e}��p���h�N���CC'�\|�r��BZ[$�H�ܡA����5S�lga>�[X}_)�7R�J�P����O��w��&!���bW\�����Xs���X��0gQ�ƙ^��/�X!��M�-�:e�؞`�v�3s�'��ER���������N1P��F��V�h�r����d=[d�V�����k��/=����*~�w�%ݨ���jB��q��[}�J7^%U��]q oQ*�/#�)���e+R�P<�P��I���f�a���-�̡-�,|zU�@�u�"���bV�ͩ��i=�`�Z��|�35�8�1,�`�a�$W��W��oi���5�mwQd |��68Q�i`���U:�;=Պ�xɚ ��Ǜk嗩�!� >�%�ŮE�nj.7�;�`%�#�B�@�����8�sz�p�Acfb�5�n�$��!��"�䘧S:F�#��=��ot�!\�XKo-�s�$�_�ʂ}D�7E�B�����/�	b��k��-*E~�
�|���i��w��&��a����~��.���` ,����w��ȱ�b�ö��%��2���¸�]�!ʙ�����+��"���;jOȺ��k�gת�D�6��Z�e��� �۰���hf(�äG��[5�Ȅ7�����䕢P�������"BI`����co��)S�s����ؔ�n���x���Q�� �=��0"�i�2c�wW�[���u�^�zwU�]�K���Q�V�A lF>�fz����B����@^Iz�CE*����aT'�u���)E��vʥ2����ؑm(��G����ln�Z�#c���b�[����L��&���s �Wa09F��N� ��R�J"���`%vf7s�>�ﾇ��W��7�z|,�X���G��#��i���J׳�fBARI�ʠ���FN��oѡ�`2�n�L �&����Q��Y�{(N�<����.��TѪ���C6��)*�\�i�uk��:Kf�=���Ƣ��Z+�nj�,pZ�u<g�C�#02R���=�!�uֹ��wm�����l�v![<���#�#Gy3'e~����̽;��*��h�{��{�+Q��6�Q��~cm��f�^+ g�!�:"�����d�GD��k5.�")�4���	&3)-���P2��@�v�K(���6�@��PX��}]Ꮦb1�?å+���+a�,$��S��R�`��В�B��@_�}�9c�6�.}yY���4��� Ŷw*gf������DY&x
*�S�
c�W���5A�U����T�R{�vi�ˌ���G/��m����.�7���^�F�47c�j�u^x̍�~�f�"�����&o�cm��L�}X"�Է��@�f)i���kL�d�W��JU�o���kF��3����f{k9w��5�a��4�?^���$��ҽ�t���fF��hFL;���[V�Y�d�I~�ծ��>��ު�}S�g#۹��m!-���kX�CA�C��~[����yP֌Du�
��g�7Oe_���7���7cv��׍���Le�H@�Ꜳ|Vs*"���'O?k®�e+
�ԊׄERX7���[	��EXE�� �i*P?ۙ$K!�n%��RjT��{�\��<���oP��r�f���
��BO"��
)��j	�o�5˶��*�Vj�F�5kX�z��-oz.����E9	Cw:ɡt��V��!������;W5�N�ۯ4��Í�[���)�ˀ-34���0���؃fQ��u�t��=c����m�#P`�Q�����ne�5!L3��V�y��ҟ�v�~�e'�k@ws�J9�ѵ~����!�?�J0�`��L�VUЂg�Z|��(�~"�g�}p�X͐>%�Ʉ�F�
Gvft^ �mCw�u�C����j� �A�ߗt���^���
����sm'�:Z��qoMV����<0c�*`R��`��ӕ�F���s}��6R�w��R1 t1o��E8RDv�P�XJ~(N����2	���.Cu׳¨S�DL\�Q�Ҙ���QT&��<�:	����"<����Z��dl���!�-OX��M[�!(U��i��Ǖ�~j��v:R�N�{P�z�V��B%qg�S�JCY��܎1����~F|[���X�I��k��3hSk�pV��v)=X�{sP*�A��F]����>y{)!(L��q��*�0���k�f�9QD� <	c�7�i9��Kǀ"�0߁ܼ�6���Pc-٠j�{:�N�H���'�ƙ��v���R*��n'Br�Hn���}�DՋ�7-������ :���^���z'�=�{���.c�44�d��0@9
G�ǯ��x��ceg2�S��'R���'�K��$H�ӠC~�W�3�s�=_NA$P4gҀ���Bj�K���?3���ŀ2L�+�N��$e����թ�_���ډ�b�^�C��K����E�3��]���8�j�͏а<.0�3��V�� �v��`�ޭ�����s��5y��56�%�6x���Y���g�$@��@tZ崹���U��y��/^-ş_w�bP~J����ϕ��=�q��8��1��� $����g�f��2��v:�X���P�s���sa��d�̓_ߌV�j�m[e����#']pA�:&��?f�eh�2eAf��'p'J��;�4 ���j64�#��=�
w��cp`�C %�I���sz0.��h� �=GgO DpU� ^��-Ήq�g2F����?�⠶��q^�m�x��O��z��;+��5C�`X��ǔT���vW��q����اϤ��LS���*|�\�o:�{���{_O�b�\��=jۑ�̪/l�0�<E#|Z!v�( �Fa}�h���Y�܈���-P�ym�(�/��6B2�5��瀀<qS[OUb$f_a(|x��?n}����]ʾ�r+Q��|+��xz�z�4��w��.C?�v�*���r��R�O����^�Կ=��sɹ�x�@0��k������3��j���+�il�&�,��k�0P��~���[�++S$�<�8���vc�?��/��<X�0��܄bR.Ԙ ���K�	f�;�k�i1p�"��i��ғL�w�s��xWj�h���e^� t� 9e�l}��Ja�v��b�������H�����)<Gm�s�!�Da)G!���k�B��DgxK����Dt��b����o��5?����D "ː#N�\�.Ӑ�Ϫ]���@ y�z������>�J���#�H ����Dc�L��{L�p���â�JZfĆgM���K��B�C����IcI����O�X%�I�"�����1�|;��Cn!�>k'@��8��xHs�
]֦�q�N&�׳�A_z�<�\���*��)�Y?�u��P�*��?;��틋�CF�g[ŕY<^�c����m���bL~��vf'�����f)ź�<Ƥ%�C�	�)A��o���n�a@���h.��A���V|g���A@^E�!���Ď�p��bQ4�졺�c�$*���ϝ�{*ٖ�(M|y�����InAm����j�_-�l�L<ba����߮�JԚ-C��*�BW��l�@��)�c�|��_���Iy� 淸_�*%�cw\7+BdW�	A#��%B'�=J@x�bK��X�����:�����Xo�D�lt==��-P(�7Q����9D��SZa0�bQ��y����f�|��B�(�S#e�FX��S���7��^�F=�Q��Ԯ�Pz]'�.b����\;j�D����X��~�:i3�M�g��]��~�K�o��Bsր~J��V��e"���qG� ���<И]�����h�����%3�I��>ԟ*+,p/�k�f~�2Ы�"�� �Փ�~t5u`{Vkb�Y��c�`@vhPP|[��T�r�T �\ؠ0��D�.w>kF<��j�2~�/�E��XQ��څL���q�>�7��Ã*�@5�j�7�NF١ǎ)��1}n���霥N���!`:*���וJ����4�� T[ =ij�F؏lyw�i"��B���<��~�ۭ13�:+�������%&�:JL��䤸�Z&�4�Z� U�竈���DU��ԒT��D�6�Q��Y���D��꿂�:�Pb{��C�"��%�m�n����ex��2���J�7�z���g2�(6�s-0H@3�)�;��llk�
E��9n�y�)W�Amcl�ۡ�¤f��]yQe�� ������?.�ґ�+\,R�WM�hv0`�oɩL��n1����?��~�X�|�2����>��#��D�7,����Z��׸/�����@X1��o
�8�S/2d'�0H>�v�7	0�?�ܾ�;,bx�B�����b�*����ӟD��6f�Fc�s��Է[�v���K��!=5b�^�pw@�-�$j��<
�:J ��#��<�h�T�'P��z�t�H����B�����x�a�����+�c��
h���9���! ^� \2�'A?�A�4ω�}���A�8���S�Z�]O�D��5Ǿ�_��7"��Q�8'�A_яn�H�c�uh��r����86k��Sr�0s���͸�;bK���<-�1M��w.TX��{Y~���*\FQ��mX��'��>� ����H/;ݟ�4V���V
��߆m��~�Y�Y�(���5����{TRW_�XNZZ�����[��tG�<���rY�aR�d@��־Ĵ[7�ʕ��wM:�z���0������{���}���:�d{�Q�N|��R���`#W��"W���K�R�{�%������$�BT;(�?�������od�WA4���"�	ôZ���I�%���[fpydAo�wi�L=]8��Vd#��+����U#i�s� t[}��n�0P<D��7�_��W[f�د�*�`����S�otu|�芏xp�oz�{n�9�V,�X��ý��kO�
L�����`�G��X���MݓKcq�+��_��f�?��^9��𣪟xs`Y+~�T�FB᪃�M)D��x&p��^Q<�e���Y����%}o��Ƅ	?��:$Y�U�P�Z��;�'�hJ�8�c�y%�"ټ� (���kȖ@������1We�$���P���x�f\=D����|#����S3+��x��4ꏉ,�1��+DڳN��SnF|�n���+�����ܜMy99+�FÝ��Z/nЮ)���0��Q�r�$�/�$�'�[۩�x�x�$Pu<����^#z�RݟSC�H�.G�zB�҉V-�^Q�uZ�fP#��m.睡���>0LӒP8HI���Z��:�v�7����F��o��)�� ^��zn���&h��]�,����h:gtE�B�����\Ǚ<�r�o���D�� ���&t&k�4�n����/����^��$b-���xʒ����^��ꡑ�B$a_ l�C��~5ǲ���=�v��Q"�NɔԸ+)T��gP�sm�>���X��I3:�\6������������{%ү;�
�B�0>a��h]�{�8]KG<{��MwvQ~+�q�͢7�Ρ�sZ
�x�n3"d��]�!_��D�b9�Oȫg��C��K͍�Mq��s�Rtr�޺E��b*�_t�.��0 ^�;$!�D\���`�On��s�w�A*f�)��|B�^3�B���v��n�.�0�'����Qd��\9h5t������Z8 ��.�����N��y�!m���g�����p�4h*`w;�8�g�nN!���ܼ4S��:$���m=J���=h6,�|c:���gø�wM8����2uxZOY�XN��4���U���W8i16u^IB����u0��}�H��9)߳��q�hD�;^�ySf�CaL!���#R�yv�Ȟ7Sa �[��pz�&�4�G�Co;ad�Lz�d����(|B�/~:O�jⰤKj��T�͈n�|�Q�����y����_i �<�������!L]�ٿ��m�14��휀r�ً���o>7�V��F|o���PG8�gR�m��7��n��bD'㤣�v�ޤ��l�z���\�(@Z�j�Ύ[�4���ڻ�] qpa���~��� OR��� �G7~��M1w���^��|�d�b��
k�Z�4�L�9���S;R/�>�	�^)x�gl�j6�  ���Y�[,	,��ڴ�/�P���β���g�g�m���?~e�9�B����3���Ʊ��<:g�X�E��%���O�wnc|��8��\y.�� `�O�g��,/�k�6�����5+�Y�@1����a�B?�L��װ�4hWXl��;�B��ś?� }K�Y��K�E��dc�u���̙�,�D�^}���>�ֲ�Q�e*�o����(y�|����̶kc��c�l#{�b�,�pQh�	xs�ʧvJ��:ɩ�K�L>�4z�ק�-��F�o|rW�M�r��$c7Ҝ�u�]3��Za�nJ/Mit[�L�Ua��:P�겙��I�)��V	�Q�����2���F��\���c)栂�`lF�)p��=�B��H��~����`�1`q��N����9v��������
v@�$��W8�Oǩ���.��a�5LY����b����2�	{��&�r���� %%/~(��38Fۨ�'wW.9tY�Y��N�H���!->~zA�V�~��M/�ع،[���[�G��-�7�-�y�:D��y����^`�P�L���+=���#���6�{�����9.�A��[�D�n6r��Ru�L����ԛ�����Œ�}hj5v%o�S ���U8��a��G�=�%�AH$�ܳ�z�~HKZ��ڝ@F�7j�ҵ��j�/#���x��2Mi$);Wt���o�~ԇ۝�c������Ѕ�˖Q������Jb#�z�I�����dȊ���M��m9�%e�@���j�Ǻ����%�)բT���ԫ}T��}hF�����Q�1IB6��B��z3ĝ0Ӌ�ZI���9�>>sz�$'`�A���%L�z�1M��l>��Ec���O��ZM��^`�׆_�>���4�R(�kUΚC������1��7���k��g���`�]A���%�t��gڡ^��l��,T�5�,2¶w�q��jfG=�ri��K(�8[��id����I%���Y�%�O>��>�聵���R^�������v�WNRQ�X�0��)��'��bW�U�?��+Mk�D�U�Z���kG���`і��&��us�����ж{n������M9�*���9_�׶�hՈϋ98�~O">����y&���Gz�m!����K
uKG���j���k�iك��X���.�́7�D�4k�ećIZ���M	�:���瀣�t
S7�\�#�3C��O�_s(�P=�Gd��d?�4��dH1�f�e�i�Γ�M� c;�J�T5aSJ�o���-J8N��q-�Z��u�!��7&��{O�k>	N����d�s�(���%�����2^��F�_�̽��Ůz�������nK�}(^��>0�5k��էz��'�_;s�r���	nϮ�}�
�7�ʚ���I�e���s6�T��ڛ���b{v�'��%<�a>�I �׸����n�5��ٵ�d���+a�`�t�s�3Ҫ���H?#�ax5�	�VN@��G�>���ɫcv����A}��5��O�Ҳ;&���P���4��y:������������ ��\	��7媑�Қ�9��(��7���*�Nl�i��E{���@O`8���[3'~�ѱ�n<�Ƶ,�Ζ��sⵙ�\KuK�j���$'xs>LN�Rk�E"ǜz�ԛ��\�N�UCɝc��..�ʇ�E3sG��}\�n�(�
��z�b��S����S�*7���I�5}�͜���n����+큘R!����
��nQ��?	������/����e��i���K���B	}9�H��c��w/%��!/��?��y������%8P/�F
�Ђ�ƛ��Zw��`W�i��O\@���&'�ho���L;���>һ��bg�[M,����*�ۜk����1ع��/=ֶ	��}75"P��W�*!�d
�!R2��%p2�������T�y�&9q�����ɷ�<�_�i�qzq��"���IH�'���zȜJ��/��Q4��|��	hi;Eo9���� =y�2��VȒdk�p�;�y tq�W�d��SQ��
_A��0ԯ�Ƭ$v�;^��i���!ݺ���ǲ�ާq��\���)<H��x�G�Y�ݼx��8��7q�c�S�#����3�X���Y��Ԟ�[0�P����ޚ��`C��#�jO䟢_���M3�J0u3�M���(u˞r9&D�<&_dw�qXrޛ|�D�}3wp��5����w�X=�S	�pV�&E� ÆA�j�}L+�cN�+"�dJ^F�� u�c�oP5t.�*� ��MW�}���:�#e@3�HbU�*���k��5c>YuOѿ{���b@�.��~�҂��F� �X�����Xs�ar�<�,�=ꖗ�+�/,���(����Ѽ��S%��	F ���cE�����m�u���>��x��I��L�����2�䇑Ho�)�P�̲�Y-�>�j�2�3^�����f�X�m碜�Q���fп�u�δ�)������M��k����:�?)���gA�r@7�g �~�%�G�c0��S �����t�}�OͮX��=,�3�τ�k��K�� ��̰�7w�tE���J�m��W����rDhaZ���ÿ5�u���
!�S����Վ7G~b�*�r�K��c�j�%��,@z�S��Q�m�	e��1�8�=��?o�ʡC.�c��8�90䝾(d�$��U���G�\���(7�<����K�y��w���X�2�L�f�L���� 
���%���L��;�:}v���,C1��k���H�2D����b�����[*HZ>�M�ʼP' �-�CE� b"��+�P�7n�\?��ü���N}~�逓�x`���П6~(�2�ڦ����ΰ�c!,z��'��.��l��	7��P�Q?#�)��Oӏ..|5
�i�J��$�t��?}d�a=�N��%�>�EhK�h����#��;k��g.���㗅����)��$��Eޔ@|6��Y=�v�;l5]E'f� SDخ����W�UK��3͂���	0��Z}�%k��D��FaE_���!�&o㭘����C6��xU�dOC�m{@S�l��`,��8�MF?�D�*o6���g��C���a�+�5��#��^�@������B2�ΰ"�퓪)��̋�d-�a�#�i���5E�<I;��'L��k�a���j���=�7e�n#�>��6���j��6�d�	}���?s�ޤ�z/��⭀��#�#�
$���M�W �ors���\2��j��t�g�/,�7Ơ�f��0�-������x0;o�/e݋�ufΏ��[b��\`})�i�ۘ<6Q�=�F�}
��	Ծ�w2�x��&mf���E �G������s�.h��v��z��1���Gۇ�����x=,�,�3��:9V-����i��A�gl:�]�s�#�K�K���s������Fv����D�ⅎ�Mo#�R<�������B_S>�T���{]��T�n.T��+7��~LTN(��D����4
v�����	j���?,b��K�l��>���γ���э /Dz3 ����C��t��:���׳dD�U��i5�����G%^5;��w��� �*;��G�l��"�ԝ�H�vl�����$8I�z��m_�Mm�5/W�U��9T�3�{�����9��>>k��!����8
͍�+'Ew4o�G�4����O%�\�f8�������#��\ԁ�u��g���Z�{8CO�H(�w�ˤМ�qEk���ȼɛs�<�y'?g�'�*�5�0;�B��9�$ڽJ��L�������v���v��I*�������u2�z �gE�Ψ�sh�St���Fb�<�����'��-�x�BX���h��>^/wOf1�P�}��V����j�{iF�6�ZFs�r�?�*�[��5�=����6,=�)=!}�O��>XD|�ȉ<�g2n���|̔� FTc(xSp=��~�mp^VƷ��X5��g��r�_w�ؖ&����H+��^���>$O�'�����媫u^j;㸎vƌ����AmEc�=��"*E�r��#���1��wmC�R M;q�>D>r��z�W�@q/A�y����{��X`A�b<��:�L�ԿaT~^:d�#�ɹzp�9�c�����׾G	�4�zт]�۟�aĭo�q5����=�|q�@s=\� V<�I�J���R�BؽD�K���Z
����F�	%Zl�l�����_�!+剏��G�>aBV��-aG��p��7�燴-�.CpH�����8�w$k���O�����d���'X��=N91�{#/ͥ��*���u���K��}k�9���"�z�r,<�����q%�����a��LVA+���n:�G���eR����d���rB�lN[�G�y	�!��M6�Th��OuŹadD��l��a4�$����e4�\����f� 1޻�RQn�Zl�
�{��"��|�!u]������T�>��=(IY>�/��2�o ��5�'�yJ�}�/�ZYd^�t$o��S���[�JW�����g��������}aC۝HtQ�s����u\���]�5 �awNo^���훽y��X3cӲc�K��d��A�+,>��~^m8$�*����˂M�N��y��*/�Zm&vy[��|j�LF�R����S��9��#mtX��i�+�����C5�6�Ξ�o����ŀ
�Z� 3���\_SAʔh�V�Ӆ\]�'݄��Gh��X���R�=$���sq���FeB�������?���m����L�F���T^�U��L6����V�����ڷ0:����K�-aO�v�-��?w���ʫ2����m����(IvH��Ե'�12EZR=qG2V����c���톒��w�ہ����N������`�Q �Z|�[�!�l��sxk��Z�Ń��5aW�2H�Qb�(�ý�XxJ�}"�+\ƞNӅu���S�<�
f���]���o1f% ���WS`�-��)�|�o�밲rV.qk~��A�ط�f��4��	��s� g�
p�j��hyp�F����ݑ\�q�?o�����R4r�f�afl�<uߪ�
X�z	y�y�N��jg�7�	�'�.�~��
p�B��>ꏇ3͌a�h�%6�?�k�姆S�}��V����*\�Ҡ�x!w�o��zX7������ P<�����~���(���'CqS����\E2��'*7�oW��g{�= ���W������\��̓(G�_P�9\#�eZ6� f�3�i�0{ ����ݟ�.,�jy<F�|;q���V��xr��ߜ͙T�w[��Rz;�����/t3��B�
�&�s#�kH}�d�>!�6?=<Pn�㮌m�Pfrx������f�Ԇ~�wo�o4�Vz	Ԙ���rX���F\���\)8p�7�TA���H�G\mM>�p�2���A��u�^��6�"x��u�I��	{��_����h�-���c���u:�!t˲���_/�������}�@q!�ԐLQV�N�W���ؾ�.^iېkab6�,	����#2ә���9�����S�\��Ȋ��Y����i6.��LT�OC7ޤ���Bq��>h��P�鷯�kR7����Z+���y+4��0/�9e������،Iݔ����^4�6�ZsO^(�S{�=7�xEȒbB�.X*���:�0m� F�Hz���q:��&﷕�˨U��� B��΁v�1B/��~��?�7������Hk�漧O>�mP�@���u�[؈3�I��?c-��0�̂�i�o�XTP�=Y��'�@��L��Q�Sۥ��Ƈ�	t�F˷�
T�Z�k�ܷ�b��0��sa�D �5�N؟6��+���ЀM���XD:1�<�ݠ�-��#�F� X��+�ʢ��Ë́���9������R��e�_	'��axM����/@�u$���G�����N$`��>6!�d�F��lk��e�̽*z�k�_����P��o��l�l��َV��D[��2�vE�)����bJq����ǚ)�B$ �wA�����N����;T��-��)U5>B5A�s��8V�A�hH8�uSd�`\��\���l�m��^������67t�g��fۗh圽Z̴�k�Ol��~���2�mQ_�S`�5�7O�R#��dly�UZ�ܡW�V-�2��CLk�cw����d�b����-0��yF��D^��*kl�_S������]VA>/�1�'/4�T\R��+���ij�<�����N��4L6Ϊ%�-�;{~Έ��L�.����鮼G�b-<6Ҳ8��_�vi�";���,TTN��bb>�E�ajJ�.?���_���^��,���k��}�4���*���i��-���{�*��<Q(a��b]�BΦ,O֟�Z�RʵS�����w���L�#������Weq�N�H�!����M�n�]Ӹ�2�,~~)�����e7tau����W��9�\g�Z:���E(��������f���~}4E�OȦ53$�������4�;b���-$��W���K����f��)3>�� ���V������#�*pg�#=2	P�.JW�&�qt�^�B�P����B}��+c��S�OI+]�^%ı&��~(��p&�f���Ƥ�E��t�?���]��'�U�)$:$R�����Q����^ݷ�W?����r�o�ʔ�z#�r5o�]�ۣN"�H��##%��:x�����]}�o���Čd����e^�5E��?-�k�����L�W�X����.M���C�Qk�X� v�����Pl_��q�#)�ml��H3C�i�eh΂���D;S2�{u�'H+t3�0?��@�
��ֆ���{�׏ � YX���������$v��~Q����	l<i}Am*f[�P��	�k#OJ���{�J�9���,�u�e��=&���[�LM��sF`��Z��f��wk:��Y"b�$�\/v���\V�?eX�
敖 _�E#/m��C�D؂;"��,� >B���rW���}hX́Z�ln�����S=���, iw�Asmk�T �_���K2��yj�Qt+�i[�YN/�s5�t�$�����!5^���X0�tǐ20�ԡ����%̲I��{n��Q%�bW�����6�s�{6Y)������\j�_m�B���ۿ�'P�+w�HH�Z���GپqF�b�i��YT�>,#�h|5�5�,�x��3�Wc��'~}c��r��w���jB+ǅ�0���:7j�	������yg@V4��>�=�ʇ��gP�aح�~6�+��~�!N})t�+�b�=���jp�,�| urM�����? dU:�gQIM�U,��3���x��7"X�?܋T�BS2m�a��[�'�Jm���߁Xj)��t4�3q���e\09M����X��QC�H z�'ʇ��]��־!�G[�ӯR�࢚p�O��jk�e���<ޛ5y�	�*|
��q!�k���c���*�4nB{yzX���F2H:��L�<p��7�|���y�ब qDd�9&7��y��������Q�5�9��f]��������\H@��*xz=�;�h$�d����c�}��[��r��͡�I���U�[L0z�F[��'N�s��Y�Y	����@Z�E��U��z�d��6�0�<K�=76ғA�m��dN:	���O��������l�|E`&���Ө(:s��$ ���`�rlꄪ�0���>�?�����˴R���A�Z<J��""}mY�{�t�h�[�����œ� �C6���E�_�����%�r�Jʙ��*)��L�݄aEQI_5k��i��l�������mB��_�C��������cE:�I����+��eZ�Gϵ�Ջ�������+h���i�@ll<L����I=>ӞK���N��ׅ��hd� Т�J����j>1��M�O������	d�4
���6B��Ӡ2���}�J5B�8�|�U�?��Ó=ZP�7�󴂗L�5 ���;�v��"�-N�R�Ru=8�e�x�t�۽\c�Q'#m��9��d��|��n����cZ>Փ�1?�+p6�v@i��A#ђ�"�!9�M>�<+�N��Ƚ]7�9���%!A�u�_.J�ͼ�5�'��@�tİ�4�e�ΰB+�ڹ);��_��O���ʛO76ab���d���X<�Z�խ��2�6>),<`�$le[����`m��Ȋ��sҁL�[;lP��+�oO�}Dی���p	a�iV�@&�ML�����R�*�:`@!
�`EFk�	v����F��$�3y����Xa�q{�A�S:�1 Ԓ��߫R�m5)���]
W������ ���?/�vI�̿�"
���2�cK����p�o�o�5ۈ7o�ќ��1�W�R�m���y(��'a�{U�!"Qq�cq6t�X��/4��l�2�w��pִ�>���������N��1X^Q|F��2�=����iF���k��MQ�;G�J`Z�&�J��|�S�ǥ{.�
�A�BWⶩWJԠ
�#FR��Ǉ��i�黂bR��R��d��q��o�!b���pY�UTN�uzdcU���Щk��:�i�#2Cu���h��Sg(z�M��p�� �E-�/����G��g�OJ2_��F�������Y����k�	g7�B&e6^�.�{X�H��r�Ew���C���d0��an�.cSl��d[#��Bw�.A{�c����`�vh$�d17��Q���'b��}��y6zB�x��|�{h�!�=]<
.�>,��[� Ce��^r��)�7Lr{cEم4M�~��I������������{���X\:ǣ�3��L�*�� �'`;i����X��L\G4�	vn�6��؆���j��$��6R���/;�/1���%�b${��������e���(��(�6�0>�E�%�����v���]�r��]���7p�U�p��_�����"��(p�����{I�JM��;=L���N���?Nvu�p�s`��X�0D�9&'y��[�Ϧ��w#�4���m�D�����B"�&�FWj�o��,�&Z���pge�x�|j@ߒ��w �p���Ij��2��9x� 9��
S�Ra��0ׇqaZ=J�]0eg�-����8�k�Z�
U����U!����g��>s*�ɼ�:4L<9�@%�5uO�����v���\�� �4��5:�w��`������+��(�ہܐ�8�"h���_��/��xu��w�yj�!g��s��YE�����bu��	[����(Yf^�TLa�l�`-W�*S��^��M�/��"u��a^3[�	��Z����H����D����9a�|L~H49?O��qA���c������I�4A=�7EV����F D����|D\�>��ӭ����)N9a��b=��$�����У�0ԏ�&[2��{�:n��˞���.[�{��;��0.��'3ww@�j���Mڲ��´�ڙ��T��T��t��(���]w5�,�3=(㖾��lJp�l� h�qQ�J)�x��u��߀�Z�
J]����-ӌ
z�c�u���`[��m���d�;��i� �}7X�����誗�IG�2G�U%��A��
���i�������Uؽ���*���b+���F-�ݾ_L6�>c�ۑ�ɧVJ�cS�J����[�]sc�Que���c2�|�t�m�v���0�dt���zg�:��Ǎ#}_p= -��a�������r��R�����)�V��}��R��B֍wj�칿'��}/�ʣ4�J�̷����	�Z����~�h?9z����9�c7��~'l��L�Š�|N���X�T��fK���W����� ���~����{v�rCu��5��2w ���R��6�S�A]��sg@
���� ��V��!��b��cF����jF0ж��%)�0Hʐ��#]!�_`F�7���F�+��{e�:>��YSue �7��ьAR��w�/f�9�A����Q�h���J.���q����.���C̞�>�:�R_�-c�5<d�(�h\��n|�:�]�ۅG;����p�6�s�Щ�s��)��g��~S��=_QW��o߻yM~�v�g�x�{�o:~=�zR5u�R���:���'m�8���o��cq~iBO��7��L���_�`��c/f����K�1�:3�e*��=�1đ7d�ǈ�-�~QOs�1V��Ś��^���c6�ď�����M�rm��{5� q|�����}$t� ���X�����"������U�r����q�6���W{Nv���up�����68'nC_�E�p���]*��6��)2��$^Rs6��+��!kX���i��4���8���8�u���b��.��wyc�wL��J0����P,p�^�E�_���u��U9�)�#�殓�*��x=!:9^I�����}����Z���~V�!�*�S�67�C&OՎ��v!9B�	D��Y6}
�����|ʋ�6�Π��G���I��2[ �-�B�X�~]��e�V�r��zk��IG��P�0I���|>x�0sW��ulgO��P�ż�L��Ɩ�?�=��K����Lf�
X��Z�|��b��m����>��(���@��}����i|���=��%�!���F�et���&IB⾡�\��'nT=g֣JO4D5hU�)'h�?,)�~�������E�G6}n�e
��q��B��=���*ߋ��ͥ��z��]s��|o-̱�?ա�P�����Q�AL�!�5��>�@�캡��Y��O[a�fp7.��̉b\}��c�����ڀ��|~-c�Hu#�_:��;�TA�;[B��V`������V�Qw��ㄈAm狫�]3b[�4�xj'[�^1(Syg�Wp���!�ؼ���z�ŉ���{���:��=���8�#�}u�L�%d�	2H�Fn�b�e6ã��Y2�:]�����{�l/�80vޮ���xR+@��S��~�k�n�seD��L�c&��>�w��S�edNNp��o��b6������C��u���Qt�b���Ĕ�#kt�mwr� ������)SU���\y�"�M�=�,�����E�3aɋl�y��l+����GWL`hZ�%`'
/^6B�yt#�N�Gd#1?7�y��#l��@�jYa�Iq�y��1Dm�"�Ê"�[t�6�n�P+p=��j�t.�>#^ߏ��p~��v��b�����'\'���S��83H��|��	&z=(f���,\�ྈ�$+{�^؆�6k�[��R��������q�D8]gemչ��EC=g�D��� ���nr�*%���+3)�� ����G`mG�b�?���rIh#eONq�QG	+���_[� Wަz]&�k��>��ab}��\�㊧�*���!Y��iE�=R_Cq�4��.���btu��t\���i�ϘC�u sA��]��؏���+]E07���:��@6���Kc�fjI�,~��k�ç���`/gX~�f�z_��)6��P�#nн��zzg��m;7�Zެs�۷`��{f[{�bsu<vе0��fp��f�ܽ�"���w����[Ä�����'�������B�p�� �\�;0�Am��/��/0��  �zG6le�1�����+I�� ���P��8�,��� ҹ[ƸD����`#���'&JϬ
��)�̡�owyvtqL������c���J70J-Ͷ \�!�"�D|�%?�R�-'HQ�� �%����|81�^����"B�:�+�~mMSXjȃ��t��Sz��Q'�bvQ�k�h?�/(��!NN��\Tú�uw�Q�g�`�$���鳰��Ԇ~+�tH����(����*	���h��G�iDw�^�I�S��{�o�T���Ͱ�O2Kr{�yYf<Z�J�O�F\��ER�s�S�<���:�sb��3�ў!%8!�1?1��!�S?��a���AJK(�T��9Ҁ�&��*��3��<���v���ľ��o}�qX�Ö��`�E[��3$�� �����Cf��b���Lڮ�$�6ŏ�0�x�PYü� ԩ����YK�ʄ��b򲬈�z���Y��YKm"���OU8d8��F�,��\L����ƽ�߅fR�V�lA�c[�"0l������$�W�4�2.DKI!���}ןN�Q8v'\��}c���9�y�}R��t�{��4 U�S�˿��#A����0����2���\v�����a"ִ8�-�����l�^ڃ�[_Fv���!��g�~�4�LT��DV?�%mz�eܷ8NT�J�7)s����ʷ�!b���7�+Q���q����'F��D�$'صQ���嫼?�QX�[�x�ZOv�#*8����z�5�CBz�|l�K�x�]O&���;ݣ��\�"c��%���o��@]��p]ݯ�`=�ڱ]�̳U����i��]�Rʭk��$;q&����m=���Rʠgv^;���_z�3Ֆ�0N�P��l�I:��.�D�`7w�	Y�8l��'��a�Y������$�S �&���f��nj�B<�D�x�n��H�ә��S�H�$����Ap���%m���5ЁG�].��HI���<���״�S���h^L�ٗed�N�s�@��y�~���Pz�����JN���ϑ�d +�?��)��OvM����)�ž��U����~1��6�W�-����~;M��q���a�D��u�;��=�g��s�B��C�Q�S��Z&��4���i�b�L�O��.+��(q��,x/M���G�Rxwܿ����>+�ӈ�(-��D�8��u���N�]q��<t�/M�[m�������ɻW�xV������#��Ħ�q�{#�����^�±	jPC��#31�x���)Ղa�P�fxӓ�X͏e]�,;B���R���*Q(Ƞ�z��k��4�߄ٌ ��&<8�@�ܔ�qܲ�k*s�麃4��.3N�����-��a%�V�(��"~����=}�i��9���t&��PH-dW���hE�MUWS�»����SI�Y�XԱ�M�icKp���4C��(b�z<-�,����[�;M�x���+�=��أK�@U�=B����kI"ѨĤ�#P�f����VG,R�g3yN�Ө}�m(b�������Z)�Ko��T����M;���@:=�sx@��4l�v��଍�����ɱ�|�0A��79��}��!N"�.�DW��3��Dh��^|�#�j�^��/n_7����rg�|`�
��nrP���*Iu�N�7j^t���������v�j�r���t�o����sLgJ�M::�����V�	��0)@���Ғ�W*`��������\��H����=EE� ��7�s�:P����)����p��lϢ/:�\�v%�U�~7�h�;o5�`(�#�>GB�Vz!�r���/K�'�*��d�y��[J�1;����[����1Q3W�����7ݐ��a M���PS�'ZEr���9Jnn��Z�3�WHCK�鎈�j}gn�8B�~���,��2��:����&7�`��m�-ߗ� �a/��y;�g�%�����R��}��dbi[�R�*#�縹X'�O��D���5�2�.X^�H��5�C��τ�^L@6�=��P`dҗ_R�F]$�n3��=��_`H������.O�j��n���=���q±���RB��|���5+[��/��(e(M-��6��NҢ�<��1��U.��#Ҝ���4�j�q���e?�R�f�T���c1hR_���쌼�lD�@����'�9|�Y֣Ǻ�=^�V1�~�����|��Ώ.���?�__�<ڥWw�U0*ڨv��C��m/.��`��\e밖$N����d �;
҃�N<���.�#е�_zJR-ts�J8t����[����.�qZ�	U�#ۢj��q�b�f���).�)�� ^�)�.w�Ù��u5�9��N�
�!P�5ꋄ��E�y� �Z�EZZ���!�Į�w^t�9��\�N�}G1��8�9R�;�c:�$�-�yMRMWƩg�jT��
��Ī�du&oՒ��ꄖ��w��Z�x]��щhJv�0�Հo�@��rT��%��iZ�;�b�er�S��}T�us.D�<Y���|X���m�q���C�V��{�2hk�啀��u}��d�=�c�Ү�Ok�L��/y�\YNic(��X0���롉��$�S�Sc*O�l� HIs�����C&���%H� e��Q�%��P\ |��J�aJ�"A����[��B��4K1֜�Q��u%B+9pf�9ę�6�7���.����������{�20��|nbH�Bj=�=���aO`�=��� @�&o
m6���(����-K&u^�
5������� ����6�R!&�v1�&cꯡ��o�n�J�=�L�'(����?�v���WG�h�gj��p �y�@����rV(,�.��Fg�q&,�3�[�^80|�����8q�#]��Jv%H��[��q5�`�ڊ`gYs�������������O6g��)��o^�%�0��d@�
�ր�f���f�j��h���� 9�V}�;)�+� �Ї=/�Q��̫ڽE1H:J��J�rq�'�X�-�-�g��n���5�F�2C2��T��6�����!��,�dt&(Uk�E��}��!�,&�+�����Tp~�}@����B(�QfM�*q=K��M�✳�՛���}+e(0�?L�u�=�ݼ����p������ �Y��������6;���Ĭ_�g����Q=`}����t���� ���s&2Y�0������=vj��L@'���iD���F�(]����S��q+3�"�)����K~����N;���)�0m��\s�0�Py���K�ܢ�d>��;�'Ҩ.H�������{��|�r�B'n"���Y�J���Q 2��0�Z%�k�5��/.�;�1�ܞ��)!j���63Ӡ��B1c�%���.�lFM��R��F��*�C����m��3���3�Wn�U~�G�,���{5r\�HE�kf�<��&������t��p����_9L�$T�Vzd�ŃSi���7~�>Y-tآ��̑�2�"�氩}ߢ�F�L�X�����'����Ϯ�y�`X�}030��ڝ�,9�)���	̢��|ϫ�P1U�@�+~?2�R�=\�{F�N�6 ��F'Iľ����uս{l�v�y�%��n�2�J�n���j)|�� �j �2�� ]5Q�� P����c&��Z�@R(_v6l�m�~���n�4�3�

��$@)�
����|L>l�����&�[���a��Ҹ)�0
�u�z Pm)J��i\0���}�D�+��Ac��<��H��5r��?@��!�!/�*�&���c7�/���L孋<�'{9�A�u{���(c�Ȅ�kϣR}�K���.���Gu���D��c�����(��h�_�h����IA�:����bK�z�ȸ��.l&,����ˡ�9N���d�вH#�[�����b�I���q��<k�?��QŁ�d��m\r�\���M���P��֩V	%yo�1��j�R����ɐ�n�/��"5+��X��%m� j�6]�/p��� ����������P"�Y���ґ��X��Y,1�ɝY`�T]"^̵��27Z��3��l��@�F8��/�����* Q�� Ȧ;�����������c�0f��35����,�7�9@���y��g�~e��&B�0�x��cL�����Y����N�)@� g�չFI�16ӻmթ���U������bcz��8��#B;�ָ`��f!
� �@97�jMVN�����هMYe=~��ل���d��]�0\���7:�m�\��� � ��h<���fO��R,ē�)^�R�s°��$�Յ��>/pY��%o��4�Yv�e&j��vҰ}��j�:���M�v�A��6�O�us)��?�B��ͨ�ú�B�HW�ښ[+E�y]_�ٸ�t�'gú��������U1p�g��T�����ߑ#!��C�.�t<�m�&Rs>�7��G��ʤ�d��pLX��t���GK�.�+�xl^G�c��������=��;TpB�|rs_�|hu�;m��M���c�9$�,3�YL�Df*�5@
��m�I�S9A�,*&y��	�xݴF�U�ޫn.�R_^�ӣ*�Z�O��R{w��sh�I��n�Ĭ������c�b%� c��m��=t�j�'C�&3����+$N���)U����^�|��/.�[��φ�~uzUywi��m��丵W�AJ'���9��2�?F?-}K�	x�*=�B�wu�{;\s:eSk��7^��T+z=-2���v�b�C�ڤ��V]־c(To�#㇅9���EI�Gț�u�� lk��nu����'y��)/���ΉX�q�3�s=/��7E=>Ȇ�r��C�Я2�YˡkG��Do�ˠ�j��%�3����;J~yhU��y�˔u�017�9s�)���j��0����+3���ɽ�]΢��3$4Χ}��=�`k�Fh#���@�i�8{����:}W�����l[@���\��	�)���E�h��� ?��\ �1L&:�Ӑf������ya�pm���2:0��T�$���̃�D���\�P�׊�lR;>�G�pZ7I�Bb��ؑ�K8��̇������d��p%ᥔ���x���X�@h�}:E���T�ǁK;�_�R�V�>׹����	�s�&��7+;g�M�Um���Ab�+�YQ�tf�KG�k0��,�m��bۀ�}j�g���lE6P��T�6í�8$��2o��`2)����QnA��}3!�Ӫ�-u�ʚ�kv�Fߛu��=o
�b�����p���q�,��s�H��U�-!���T6��D��9����&�2�7�1��C��SЄ��A�����$S^��vfMz�Ǯ�_�^����������)?QD �yI��ɠ܍r溩�~�V׭���<u!kή}	��I�f)���x'LU��t��<<������P���K�zs�����3R�Z�
�wl���7��XE������&��3�̇ӗ ���O㯀PdX��EV�RD*>��hp#i�=�*8I�4��
C\n��Bn�Ѐ�#Pv���-��}W ���m���;q�v������ֱ�r��ah�\����)�^q�7��W�J��>4˦��;Q��-re���ܟ�hi[.�蔣��I_Z��Y!+�n������[[�6�v�������)�&i"��a ^��D���*�-)v3�	��B���&��H���}F!�o��H���r���4f�k�eRj�j����I�&m%�j��7:�~�H�un�Od	��NĂ���������WH�/�Bʹki�����։�.�1l�i��%�Cx1��]��x��_][䪒c���D*�͹�f�+ʴ?'��:0ߺ��	�G������:�g
�Lb�V�D�8!)�md�ax�^L{T"���,�uH�7��^~����|�Ћ>1��\s/T��[L�D��.jQB��Ik���tY����X]��9�߰7���NB�/���򦹴�7�B��.t�Z=_	���V{XH+4>��"���r5����\I0d����$�lY�x��uN��b�>�ol@�Ҹ۳�U�|o▁�G�Gr1����g�*ؒ�<��qAQ3��)�,�$�DM��%!��m�nP��a�l�]�K�Nk*w�km��5�р (*�U5�4!?������`:���ɺ�z���9��'�����X��3W�쵉a�HǛL�d��:+��Rؐ�(��ik���_��Ùrp$�Ҕ���jA:|A\���J��&��t\X��T1a���!�
����,��#�z2��LV�đ��Q��fIsJc�V+A�����L�˿�i��<<-��;�N[�q)��G�7�$nSX��a���n��g%F[�]M)Sr�W7[KX���:�>� &����K��y�jU0�WX��^Y���N�zC���������҂�A�:�I��<�FX�{��9��Ѿ��T���kC��$F�|\%�4t��@;I)pJD��lVJ�P���Hp�¸#�ў]�m�Z�:d��ϐ�g����:�u��8/�����l�7�e��-���W��5@��=�a�:�ڈX�-k�u��{���$&����E�[�*kp�6��މ�x�MQJ +t���r��)F<_�:�rAu��DM#�qQ){;��W{���JF��NfF&ګK;�y�D�C��5dR_.Io]|�4�S��arM���C莰��AT����M��%�-.Y�����lR3	e-�f��D=�;���̹�m>	�~�«�~�%>sj�N4�>F!�����8]\2�~Mv��n\KR���󓦷�	������l���>x�b�
����=��\Q�pՃ��c�_w?i���G F~S*��iP�+�p�kt�٪O�*t�����z�7d�P�;�������!�y����Pc�^�+�k�:#�!�C&\�ϼq;J׃�(����D���}%�=�:A� DT<a�1~�tXߔw�Џ����1j ��-���Ĝ�fJˠ�Q+�چ�)a�-��S��s�[���--��H.��G��v�:UȜ�$���F���a&���	rBT��;�_*�LiKY�Qq���z�����ne�fitM�)�1	o.�L���V����b~T{�M5�o�Q7�J��Nt�U$_6Tay�۰�]�k@q�����/U���`8�]�?3���M�4\Wq��ћ+ݽq���T�g� v~��y$*���qCw��aB�km^����~���ϸ�x�B�(n>!XwV�6�ɑ�>
dT�/8
�=���!R}��1</�Va#g�P9e��@�u�{-i{�O�P��!N��� �� ����̭���V(�5;_�PC��7	�4����A�u~�R`躛M�q��\��N�s��t�c��{9��
dZ��Q���i����5]�@{�0'��-�g��\�^������=[��j��	8`��ףCdC��&��'��t)'z)�5������ay`����)��"d�!B�z�p�(��3v;0luJ&����`twZ�2ޣF;W��U�~~�z�o�N��!��S�����b:��k������ky#�g��3���D���\�}��Z��鶸}�]u�F���'��QU$*Բm�B�:4������a�����Hn�S�hq��YP�Ɗ����H������N�,$�0�����嫖�;@"͢0EPi]n��`�i�w�]� ������5�dwk�0��^Ϡ���([��=.���h��B�Ʊ��g�h��JA�D���P�;�֣�˶4�e
�ށ�C�xly���
]��1���V\��Ѹ�ԧ?'����q�z�i$
��(�h���69�.d������k�X�{j�.��VC#ґ!~�T?jԠ�x|��I"q&��pS�|j�l��l����d<�8h��F3E[�@�uآ�Ym�i� FB������L.P������JC�d1��mm΀�����r44�?8OA�&���Y��8�~��h�w���DY{�m'A��Cz.ޙ�D��&�Bn�����g�����q�:�,M V,'�Rٓ�f��D��M�lT8M����r�(߆8XK�3|��wZg�&���au����M�`�^���Ŧ�Zx''V��I���r�ɣ/��F7u�}m�)7w}D2��.���
0�!� �N��%�TU�:��6��*<B�L&��l;8��#('�m�"�KC�&�����oX�|�����e,P����)t��=mi����o�K����"�뱐 d}���`����q%�����)�4�cb�&��W1�s��)�2�f����$m**!��B��,�nk�ը9[��wL}�x��>c��H��v4`(st�e��!q΢.!�Fb���O�<$W>�m��
��L�2� _��C#�}pA�0�_�X�K�6wvz��:"%�L�@$��&VǷ�tQ@.`'��7ܼ�~��v�F��"�����vUzц�g�!���<�����r�]��]C�&�Cb����ث:���N�N6��Ç=^	��.�)/�����En�HM}����S"�VZd�[Y'�����.=ϸ�D�щ*c�J�2yU�uE*�@	�T�~���a��ɠ��g��Ԫ6�
gVX�[b��VC�2:E�'Zق��`T�4�{AX�4��'6���-G.���{���n?��U�� ���_nm ^�$V��%��Q�ϓ�z�B��z՞����F�RA=�i<i�A����2UEށC�5C ����I3`��	6\��D��D��4��,���#��l1�C�>�I!���O��Oa�dݎȠj�Ը���x��B#-�W���<P1*�U '���=�����L̮��C��ue�Ũ�Ǣ~��謷�J�x�٥�*�"A^oVe���w���@��٦������J�xH8�V���|/��W�,�0>�J����tJ2G�j���Wb�4����X�ߛm��_���|�1�d�>�M���p�����U6���VZ����1�|��l{�)S8�rQ��4Z-���'����sIw��M	k�q悙쾸T�{�� ��W�b���I�,?	2��kᣖ�4�N�]F�W� �E�����ت_�V���{P�0�m��Ļ�U��@:�1�r����aRU��n�B�vc�;HPd�M'��ϴH���w,��k�b��6�䠖v}8�ȿŧh�{����0�a�2~��T_���g	_f�z�kb<V������eލ�hz���@�,��m�|Գ���5Aj�C������:�t󏿭�;��8���]��������c��bm[��A!�M`����DhA8��'Ya� WmںFmg��������<��qe�Ɣ���.�c��:xW���{��c	�֭.W�ҙ����I>�]����%s�Q�6�J����&B�u=����&7]��L��<�Z%��;X3=X��G��=s�C[�e��j����	�|�D5Q.?fS�9`�;}����Ї]�l3�/��-����lrU�|� m���0a���"C�7���\ͮ�����:��g~	�G��u���w�����p2g�Z�`>��=�Q2N����<X��󀿜��=Yf��x#r�b[��X_�C����S' *�P���>@I�J��p��1��`U�k6 Kg��mQ��ТK����R��,2�|�ruQ���H���o�;�|�w�*o\���p�)lL1L�(�E��[�d1\����q��^>�!0��\Mt��o���`b��>��k���9,��T�-����=�1+~���s���D-e��ϔbF>1� ��X�>[�_}�9:mͣ�X�Ֆ-QW`M7Qj�K9m�{@��r�drGf�J���I��Z�Xt�Ǟ��m�&�z��ލ�8����<��CK�(��~A��Tg���\��#Y�ň���xIa���5ԷSO���G��D��_�+���`�tw3�=�C�(h�s�#1 eX���r+^K��A���ˣ�c��Z�ԧ�rIFrA�S(��&���oUi����n0���,{ǝ�M0n+��G��L����S����/�]������m 3̉:�S�6�:�䯰�`�<M ��lG�5e�N��}��Ɋg� ��cNgjN�8�jky*����a~@�0��bN���O��:@�����D2�2K��� +�G�E�H��\F��C.�A%�..R��� #,4Җڵ�Ϥѯ#[i�|�8MN��~��\&[3r�����/{:�LѢ�X�qֹbIqv0��b	{H�OhCXŸ�zʅ��<7弒�r�/4�(�3f�@S��h@i 0 D�f��'=�������4����Ym��߬1��* ��/����pGFS���B�(��$^��i�ZNzeV�nȳ��F}9��q��P:*�D7��C�d��OM���\5	����N�ȤX�+���"@�r�p�w����Å&
s)(�����<&�����]������>?�yn}��UY07���> �&�����L�g�F��NM��FZ��n��4J�L~3�0Iؙa�!R����3ѮyV<�[�F�W�Cy��`\�������N}?l�T�|]��tDO��rc7RY��
�8�[�|q�g��U��7($��D��������rV�4��m�.l)��0���}�U�����/:�>2ca]�YqS��J�u&��e-Il��Mo����B��(.�{(�Sq�ŨK��"Piy���&�+b�ܭ�Y����l�r�A��=����W{�̏�S@>H�RȨ��څ��I�O�yRr+�/�J�(����&�;U$�֤��ː���=Ȍ����p@������bS8�d�Z���q�q��wz�43�a9ͥ')d�nlG�܇�1��W fӥ$�����hbA�9Q��y��S�5���Gq�Fl犴((07���������ht�>\���VQ�"�$t�Հ��mlޣ$C��i.����.~��-�A�@��L�p5���!5A�U/Ǎ�Y-�;�R�����5��T�ƅ�*S���?����d�2��t�?M�L���p��M�I�ܧ��G�P~�4��7pW�xp;*{�@�E�S+#k�m�rԼ2��Q��:��Q:�Uj�tM��$H؁����M<b3|�A�� >�B�ꍦ������c��YzQ����A���(���W�Haؙ�16x�	zI
�x��<����y���*0�����F���=�>	�l��x�#��-_�_���*�#��)�㚎���H��A�8��E�
�ԥ�d�}�	��.*B��:��=�v������'n���;4�z�%FA ���+ʪ����ӌ�����2%�[/P�8�K���<�!��C�L��:��R�����b}���o�q�?�=ʏC������lЬ��s���e4^`֚s]��X�9�M��meqq>a������(��#�JaR7��G�Ci�:w�-�w���? ��8Ӂ�kJ4��θi*z؁��.�A$	"�[�Ja)�F���g��4Vy���,
Լ�k�2�3aU��j���Ek��GCs�Uk ��J�z;C�r'�����S�����.��I	�Pg�e�;L���4��V+F���*����Z����?G������{�l �D�}���k�gz�d���9�й�x���_G��a	��ǍX�B��%���Y�!<����
�\���w�č�p��pne�u�J+��'������d8�1��Ô�H֭�.�*>�=��� �ɟ0���!����{VU��s�9��@L��ɽ����$�dU�~��4��Zə�o3'x�,Fy�m](���ՀB�	y�B���Ѽ��*7��͓ȣ*"NJ%o�gM�r3=���'W�M�|4i���r�?'-��H��<A�<	�ǘ�C���9�!ʂ��2-�[b�� �r>�G��F��4*�s��q`���������xT�R��UP�c�䰕v_�
1P(�R��.����G��G���d��J����\��._���B�g�h
ű6���f\<��1�7��I������b�bG�φ�Y�ٶ�խGJ���T��VE��Y�OV�=�a&�>2l|ҿMo�r��7M�XR����Q(bX}�R8�M���y�8�Qξa�9��֕���?�#�H�~Z<���U����H�w�oR�ϯ��}LjQ*G�����~s;dxDJ�J o�*l� a���	�-CH7։6 =��N�:�NS�Q��9����\�&��FvV��M��~�ǎ�Wu���S۔�hѣ}ߑ��)��o!*���z�����_ ��.��ch��Q2Átw��4����J�=�RJ�gW	T(��`Pj���n������_%�G���P�����PWc����������$���h�:ߪv�J��v�N���Z�`n�Y�Ё��*���橾�j7$'&�*2!��7��Q�ƭṫ���F�S3u�����4����`d��<�|#kЯP�����o#�DJ�i�w��H��f��ϐ�����{σx�A1&Ğ�0ӯ$%Bt���:v�M%�Ϭg-���K�q�
o����Dro�W�1�.Efn9q�1��6KL�x�FyڽUjn�[F��=v�>�\{@�E��c�G�;�O\P&o�^���Č3,LE�%«���G�U\�g5�[:�tĒsWN���'�|���M&�&Š#�Q����<$zⴊ4��ᤆ!OG�mXs��������
C�S�8`�0��߅��A� ���nZ����@�_gﰟW�h!V�n��� ]?k]���ƌp��5@ �6��iF�lUޘ���3]� ||�Y�-'�>2�?$g�B)�a�����.�X����Jp�3�M���r2�Y-=h?9o�k�f!x��A�=�������l�"̌����E;�HD>hR�p��"�OA��i�3Y��3?�w¿�`��8���j�Z���b&<�s�m������0��KM�ĕ�M�b���ã�N���7,y��z��9�})���a+�Qs������s��v�>��Y��k�x�FRҝ֜�D3+�_\dB��U����R&�r4kV�6м �d�d���՜\�"�s3@_X�a��0�zy��u78�I�RUF�94�Ie}P��k�R_��,�n�V7}�]x�+>�M���!ڥM|edT��;Ҵ_2��ɬ���<�XFG�5 �l7�xaO��V�\�M�X3��P�;;	N�m8��+5_��@�2nܲ� Z��4GZ��>^Å������\�w�:��'��_g��O��!gp�b:������
�]~[����.�D�2����GN��
���^J�A��s���$x%�]a.��)�b��![?U�^r�����_�ZW$���?���ռ�B,��KU�;�6+J��4��2~�4���	 -x6��*��}EK�t�k�:�I"M#�Xض)ϣ��������*M�	u8u����� _^Ng����]/>��D�"_���mo�COl\1�H�����A����Mll����`�\JnK-#���K�H�8G�ʖ��^������
5��}�F��W��e�ܖ��ϐ�2:y��戌aO�6�A��A��K�H��1�K�>O#����aj7�� 9����x<��X<�|N��v�����l�`���J�2G	/ %��e91"f?��A9r�����#{��(us!!��-��&G�Ȝ�;�Mte��z���-_W�QHG�̽�q��T�����k�f��S<|b-Y�:�Az�,�l��^�+b�Y�4�E7G&����y�ߧ)�Tp�۱Z"����������m�\ˍ�#�n,漆�7m2�gtAۺ��US�
�y��/�+���^�����`1�!?�Ƽ�*^af|?�"���IM).�=lfc�.���%�+����C�)���C��R�[#��!Q^� �h�h*���ɹH5�*�S&�.(	�����>Y��x����et`�R�S���4tRa�Q�I���Q/s�
6����d���4\J��GH�Q��8��Λ��]C%�m�%��n�;3zk��k�m^��n��]�"7�K��*�Cd$�{Z��Ő�����������p>XkT�U�|ʬ�.3<�e�K�d��S=(c3��+�筆۠���vNS���s���v���-�E�;ɴ	�=|al�6#��eb)N6��`������۠�8�Y�_%B'z�rE"�oC�	?g��:y�bi����^s\�9�럼Uܟ�lͅC�8�^a���}�Yd�р���9�;]l�D����s�
]��R	��(Tr
iPZ=V�l��/�sl2t�u�[�8f����=�qEul����d;��G�=<�F����]�9hae��H}���r=PP�Z)K�9���hU���L�=K�ȁ#0�u��DM�`�dˈ����]��ȇ6N�I���!�1I�+T��i[��l�>gf#P+��=H�ť�/���H�j*0�E�*dQ럖3z���Sv�b��2E�׭ݟJ���ͅ�[�f �������	�*�H�L���˶mM�&q�<��]|�=���1dG]��%&�o�}�7t�}��v�n�
޽���jG�T����/��L���G������둂�O���-�:�z_ �ɱ9�<[����B���W;֢hொU����m�W�i�>a�ym4#��w�Qq��e�~k6"���d��	+)�M���'���@�v�Cp30U�E�\M"�R?�N7ϻ�|�P�^Q,O���z���L3��:��f�ڈ�;�2x��>�Ld�҆��_��Ĩɝ;�K������"ݰ�]��+uJ`��|�����V�ྠ,�d��*}z�����~���L�%�bM�CW��F��̲�J9l��dr�2jc./�ӂ;�S�\�D�U�ErT03X�y�L�Z��T3��]P:?C������+f��7K����͌j���P��<��r_��B���HT#;�����>��Q���rr��zVX�F���8~m K�a�E>�!���!��*�P@��&	3-�L�#6}S��>�ʾ�g�k���i��`.[y��Qda�֩!EJCPi�ff>fF��ϣ�z��ey��W��(-����XT�e���q�-��D?�ڗ�N�e��Z8�q�G��|��J"�å�Ǒ���,tu�J�ܫ��V�^p��p��8�.a���ĕ�c��;B�,2����v ����ՌPh���\*�V ��-��:���X����~�1:�
w�����E�0�p�w���B�����å��
�g����I�*}��"0)��7�7����g9hXö�*��=r+�Uk�t�e�(��8�7��-p�[#c�;w򭥘�m�wv�W�INO"�Ln��U���vFʣ��98��8�9��Ԛ:k�'�� Ϲ�h�o�����%o�Fp���I�/!7�z��v��C`=?:����J��Fb�<���J�U������w���� �{�{M�4Q�������2�P���̪��T>k��f/k��ޟ��>m"���5��ɑ���;���,v+���QԾs�B��XLv8��<�zu�E���^x�t�C�)�\o���6�~��e�?��e?�8�4�z�� r��1�Q����!����U4�f� � �0�rђ�jө�`���2x�b����X�x�-�BM�;����?$��a�5����r},a����r��I4����Υ���)�E�\Bђ�����<�AOu�8�G���ȍ��G��2���|�6��B����Y{�<E2��CZ<�HH��������jC���@��b��J��V���+Q��Y���}YZ"Qy =&��\�	�tR������l���$���l��6����>��Z�Vݳ_�:h�v�
u���R��y�u<"'vz>�ïb �f���V�����}Y�����aHR=�9�SM��tG{|�8�XX�䎲�oF��>���D�Z��[�2��T}�M�_B�| �"fKw	��R�*��ߗ�$���WE\�=��V0ke�6�d��Ѯ���ʹ`ך�-�g{N����{�쨛kZ(5��r�[®��I#�4�Mth����'�p/���NC|du��7$<�%F��vK�#&��a�cF�a8;����^f�2����]�W��7MJ�н|ń������8�Jy�Հ8�W��30[|�	4鶦4���~�T� ����m�(�(D)�2|�����287e
W�<��rciFx�Yk��~K �R/c=E�q�Ylle�,������jq�9��ԟ8fUXY���u"�E���0�Â$�������i-xYt^'�\vL��@iq��HuR:�� �dكJ<qs�2���O �̷�y�jD�MY)@���`(�$2�FR�!QGl_
b �A�P�Z���w�h�Vڞ���<_�{�i훽��_�$��6�!>�mq��	b�rkIU���B�Ӫ���q�<كw��?X,/l���X�����H����E�=���%����I�c�v%�`�;d$�s�@A�q�xp����-�,{����f����8n\�=Bi�
�C��ܩ�Q��s�Cď�p�l�VE	����|Bt�7����N*N��9��kR?��<J�|�FڽPCA/��^dq�TNʦO�a �<�}e�tm!��d�.Oփ=��H�v(0B��H��w�>�x
ZC�mZ=5L��o;��� ���>
�b{�W� ��f��R���&�B��l|�m�.wHn�$5�ڀʬ88��Ǳj�h�&^ɠ>'q
�`�:�X9�$舁��&c.^��3x��{r��#pݫ�ozs$,x���G��~����U���'��e/���߂�-���(�"�Ѩ.��ax�G�og����
�7�r�d�D�������`N���|.�D����MlZ�h����_����R85�}�5y�[AT��D�E�}
i\0?m� ��-`$]�[�u��V�1���}7K�5��b�q�[���<��_�/����~+��&���z�kq��N���c��[@��į�`
��m텍��'�e�Q̈́�ɷAvﵮ������b�6�e���{aO��q�׺Q�As�*8l|B�ۧ'�D�b�P+���*�H>��X��n�p���h���'��fQ������Pl&�!�ڨ��d\�W�F�F���$ez��S��:�����6nIw�5꠮��|Z�V.BN��?wLCU� 0ϢKgE�#�~Y���>Ys��eZr�3k.`�g�*%P�P+��k���V.�E�➝/�,uFy n��7��Vi4��z�!dK�-�	����>����S��d4��[�Z���G9e.���CTw>2s�����'��ھi����F�{'��[�`0��������,�~ҝ�S�S��&�;"�m��|��Q�������p�x�J���B��X=���_5��3]K
'4I��0`.𮛃�s�m�����e����Df����i�0A��.1���\��§�)	�օ�O�LN���A��D�� ��qV��ZT�F�`f|�O�ȽO� �4�k dޟԅ3X��#oW�'�%�M1%��O*�����>����>4"&3�a�?o�3^ܞ�,$=��Xz���k̾�Δ2�	����Rή�"�'�M�� ���9�"�>j93���6��0�d�S}g�SM����r�K��"��,�w�E��N8q����TI�S�\/�jN�����n톝n}�#�tdl�`�H����XT��d�&��R�XV�I�����7E��*�C�m�������
�6!&%��l�(�m�H�C�}ް���h���;�U��@�9�ƒԖ�#*�x�q�
�D7�M΅dρ��]��)�&#�dz������)|�c�0�z�
�ƚT��������F@f�K�Y�d�i��ǹ$���Xyt'��2�qbD�ϳA�w'.�?6��jM��JPŔ�͛��dh����׏.���¤�ޘ@���S�_���l�і��{؞9���j�h.FIz��p������M��MP�`r�j��Z���o�|ֶQ��C,��B�Aʏ�ˁ��Fr)T��J�B��K��:��5	�,�`k=MS��	����A
J�	���$����G��r�$����?D_IA4K ZA^��b�;���(�@an����8���uB��Y�xk�lߠd��l���ij���5�c��޸vL�툊��N�l�ܝW�;yzDt�6}8m��~��*Q���37�gPk-�VqO�(�Fk�8��a��(]�3_ߚ�[�J�/sf8}�d�{�N�bzk]+(i��p��X�����H��>a��/R��Y&7s����aYO������Z#&��Ãr�`�C���{-"aAH�2(C�������?����<T�ԒQ0�X�(H��#*�	.ymwX�'�:��(���~�Ō{�}�56ؚ����^��x�&�C��6I��R�T�u=����IQy	x�n�qwa��p��;[W
��R#���~�_Z1e��O��Sv
^�tw0ΜX��{���[���U��E�A�7�0L�nN<D�)�Rfq6��;Bia�팯W`�ut����n$08ŵW�q�^=�:�x�M�1�Kl�1mE�Tw[�vL��Q"��XQ�2��Kq��N��z���&@�Z݆����H�İ0�u���":Obk�kW*0s��V���vGl�����K�.:����y8\ڛ/9��ICh(4��)2ި� ����i	&���f@<C���Lx?�ŏտ�{���Z��谨�"�s&$�ۅI�J#]T֪���oW8W�Y�������n~2u��=RL��m)��VCՠ�k�'��9����j��C�i���yB�]-���İ=U��r��_�q%��H*I�ݍ {��|�� ��_�C�I8r���C껺�=Eo#N-���;ٝ��S�Z�蝴�.g��O��t�"��|*B9b=�MQ��#%�� ��}]�xF�PT��ն�b���Y%5�9;\�twX'3��b�j�`)���3R�B��;R���=��7�������$� �_q��DG�ڒ�E}%J��؊�9�=F��K_B���IE%��3��������ZP�L�'�X��.�I�U�z��|��DP��8G6vR�	>���S�L�s�pm��1�n��|m2�]�F4���L�ұ4��:|�fo��C�}��#�;�-Y��^
����&��<s+u
�cĶ츒��)�H�\?IW�pe���m|�UE`#t�v���ƀ�F�K���Y9O*��5հT!��-�Nґ�k�}�x��� D��H>�����0�Za��|#=;�r ��r��>Hw��Ʀ7×@�&��`�2ۣP�3�&�C_o �_�(|	��K?��=V2�E�RF#�w#���GM�����cC����s�|ջg�ȑ&A�Ԕ�d!o9����%D��ia9��B/!b䒸�A������y��Gx���H&d#�q��ludQŎҴ��!֛<�)�ڸdB2����kxGM������ ��@m����U�Bx��Vg#���|�(��"���&�m˭��5R��2�'�%n�i�~uR���X=�a2aw�u|��l�\<�WUE5�)o^$��F��N�6x�-��bU��8��7&�:Ԡ��=�D��(yI֠�wb��mު�u��r�;��:�|���:�P���M%�^="��8'���,7�8�����wNw���L��&��$3y�K��~o',	��'��z>�B�7�8���o)3�ͧG�I��'1>u'k~�+��X��	�:إ=�� �l���S���"���,	n�xi�ȼ�ԯ/�#
i��6*��dX*�qW�L��Ƭ�;��Pd�Y|�2�}���5@�U���>������ďmrU�����PqVM����Avآ��^������\@��YD��i�(��Ž���șz�iw�B:l���R\�	fo�"n}Ŷz#��~��A���Ơ��g�G/�@�S�B�@L�_�CN���(��޼?2Y}��*E/�90D}.�A~��D.�N�lġo�x֫�I&���6
����8f�%���iI]��������e��A�nV�4������k��Fܽ� _ͰsϺ�/�Zr�h�	���Q�A,iG�V������ �R$(�C���?6��W��$�Fһ��>�P}뒫��A��晙6���H��8am� �	�o�rzc���>U����A�y�Vߎ!X�L[[Q���|�h�������dluuHk�n�Uv�,t��TE�Aܨ�ޒ7�F^Q�#��\'�E�C�2q�-I���VԌRI���0S�l-�Bk}~��t�92f��>���cG�x�5gtm��C�B�[H͑��'�((	G�V����}��P�
^��Wa��X�J<DQ�
�Q�dƭ��>�7ʃ�3����ß�
�|�f����T��5�ۘw|t�xg!��p�m3�g��U���bʈ?���>J%�P |=a˛�Lgn|�:�&����VI�7����ʓ�<�͵��q�Ѿ�-�ڴ��e���|�3o.ǹK7���S,0/j��3@��}�\O6�+�>����*V�Rl��BCu���
ʜ
@g�*Zn����HCh�@�Ԙ$J���x����p�Ŧ�� 1��`H{���������/퓗$]J����b
��6ҟgd�;��wb�F
!�����K�Ol1m�{��
͆���mu����Y�1t	�Q|�x��#*`QZx[ H&\�n�?3�԰A��-����8�C5F�"��5y�m�E�k�) ��"?YZC��>�����d�6|����j6��g
�y��3^�������7���d�~y3��� Y\��^��'U��g{/2X���6�j�����\8g-C8����v	���~�cr��J��<D���N���E��]��kq2�i j�:\��>�ex�s�,��1p�7�m����p�PB���u�����d3��o��=D���㯓G'Nn�ˠ����D.�h���1xJ�G�.ew�����Ã^S�u�����,EHf��녚������G�K������`-��W��U���'�A ���<��������9��e�N�a�X�a*KbG�eV��2��o����Wlw�U�q�������&�E�K������^���I��T��T�����a&k��1�e�?�%�ʖ�vM,;�k�Jskn����j��r������%�Jij�%#��vp.�U}q��3�HTm?x�����u4�	���q��+[s-	���� ςl�����`:S��JJIy�gՄX�1�b�zQк�#���9�j��7R;���X�{��x�s��.7�T�ߴy�kR*]̀N�k!�����u?��a��p|���xV4��Z��|!�{n�#b2�JU�	���8�qb���@��T��-��9V��=����_v�?�̞��ctL���4۬�.W������u
���uqD�B�J4m��E��P�1�W�D�T����T���H��л�!1 ����@��yo�4 մ%��r��R���	�`,Ҷ��\1X��D�a_�����z�Ec����MҐ�o���*Gix����3�J�\4�>n�k=0禗/[q���|���#�l��K���A|-NO%�M}���i_��f���I��|�`����	C�c�� &zʒ1���y ���D�
�"�jn<Gg�s^J�$��eDa�fu��ܛ�#�s�Άi}�f�]8A�~�ws��J�뙿���O��7�P.��βz'lѷ��"�*��+��ȅV�: _�j�����3����\���iG)%���X%����w��Ŝ�E�.
W����年��~���_�eH�N?���������Pab�gdڶ���mqq	nh ���8����$����K�ìW;7W�cl�=��h����GK@�-z*3@5-���z�E"�o�낰5�������1����WY�o>Wdau$K�x����
�aH�����Dzl��v�QdV�+ɪ�(��c������e�1�GIU�e#�7?�~xď���;�P�秩F9�\�&����y�!����[��n�Ra�3�,
��-���-0�� ��f?������dðjc�z/��Yd\&��g��huݞ��:DVI��؍��Sx��B+�JY��!F_��5s�p�;��@���+�k����?T20�eIoHz+�S�svMb`���	�@�Mmy&�2�x1�1/���A��G�OfnH���0�V[P�u��ʕ��4^tH��^���J����ڝl�pq�@W��܌c�q���k�-�z͐�L�o4 )ႺC]ɡ�F1Cwr�p>�z ,i�s��[�����/���o7�>��%�,'��D� e�����`��S�Ҝ�Y@�i*���T	]�����	4᥾}��BY뀛�~��61y�/b9���F)�j�e}��y�iH���5]�9�(}�uk�ײ�\��8y����
������p�����c��p���:ԕv���ISI�{ɣ��IQ�g='c(Z)	ലd��0m���(�;�W0����5�9���ܞ��4ءwq���RK��ֺ���>v�RԒ�T+#�G)��2k�O���-�Ɂ=�A�nH�՝�1Z��ыO�躂�:/ a�:��5V2<Y�c��7�H���Bhg�S~�޷}�
�J�s*���q�����nTjl���E�gҋz�vO`ҁǏi����d���o�ѡ` ����ع��s!��u���N��ؘtNV��x�	�9�!��s��}�:	�?���ل��2�q�uCUո?X7��-r>�-�4��N	P�p�D��Vb����J����Śc;�$�+�Xm��6�����^UɶA��oDI� �|�a>}���>����j?�8�>��4u��$sz6�`�v���,����7j#W���u�n1�����L��������keU8���P؎$��a�j������E;(��P�5�z0-��[��1�8\��6����5����t�7�l��^��ِ��'V�SwMYJ�
�m��"�]]�R�R�~�W������I����3k����"�5��UZ��g�K`L��6��g3u�l]vK~'�|�hǲK��O�A�1WP��d��H��Y�c����|(O���U���.Q��aD2��\����89��X
�ת	�<d|�k��[I)�(�9]=�n�j�s���|8��S໇K�@PRF�.�(Tn���=˟���T<��04�gn.�X���W|T.x��c
/G�O�*٢�|D	�2��<d,�{���g�7��^/HR�#�H�?�e��nO��Zc7'Ԝ�_��C�e�{$Xw%/N~ko�
���#^5������L�������
��m��� ў�l���Ϩ2�:BK����� �xsH4����7�r\�҈a�8�W�R��z�� ����HH$sm7Q��֖iu2�V��Qpm�3 ���ś�`^�K��3i\\� �tv*t bfz�Ae��J�~K�۵�g��݀ZB	g����\�l	��okZ��	�� e�?98����Y���O5rh�9��S&���Js���>�?��*�3^ (	����t��p�̜�B�?'�Z�����G�ˍo����K���j>!��y��2ٱ�Vsn��r}�q'&x}.;2���l��'�~}���VG���ѳ"�w���a3����)��UC�a^$>d��{�;�ud��l����&�@A���'!w&���o��WF׹2���w���]|"��Z��s�����z���m5fh{���Td7t�o�D�_�*0��üe�=*x��d�~ŝ�R�s�`��	��*am4�e�W�]��ˠ99o�}}���f 3�yȼ�6,�:�Pc`*\H�ş����W����m�A��>e�̼fb��պ��ZH
�0[#-�k���G���qu�lط4���W�R��\k�u<役�&��c�d��D�^	�F��w�gE�a#�?�蚰��EA�Z�ObI�-�:N�$�zJل��ig68�`��n�Y�!��:�9��]���B�Ĭ �As���������!1{)DX1����uB�2��/��#{Ev�/������5�f	Sa�VV��c��IF�]�s~�!�ukG����OxH	e��e�j�^jnҎ/�cf����nd[�ov�NؒSg����`z�w��k�v�,���g���R:�ۂ�<���fUf�69�q��)���^����������pF��d7�)%����b,��l���4u���,��>)��AL�W���O�@r`-��:򤍸>��ķ�c�[W{u�$�Mn������$�@�0��}���Տ�,X�-�Yv����/�#��%�j�edS-G��'1�2�ܙOUƴ�p��##���0�ܖ$�S������8Z�>c���$uX�+���"�����T������?Cze���6�B�=S�CVK[u/$�M�I�9Irt2�����d߂�:e��%s\�������t�p$EOD��N���c2=�U�'m�rT�C�F۷g r����~t�ً�A'���H���LКc��S�)5���
�����k
$�'��b��|���i�Sa���:�N�y\�����M����:�:,����hZD��Rj������4�@�(���x�i��ˏ6Z$;�hSb\���M����K����J�-��	�O��g_lI��<ׂ[�0���G�*���B.�X������)a�vQ,L�y*���}��&�X�������b�r��]�=�7L���HM4��p8"TɊFW�|�:C1��ZHՃ�ςE�pU��v��*ER��Joh�6���V-�y�$g�&��*r
��s9e6y7zp�
��2����'sL
�qSs�7A<���wAk�D}��c���t���������-�D��_��W����({$��LsC�v��.��J��� �����^iڋ��⮍/d���(��ffQ<��&n�m���F�߈`��|�P��4�s�6ONx�a����$ $��VɃ/J�	v�|��6n�B���L((�V�i����T����k5-B�hƗ%h3��~�eR��5=2t��$�^��?����o���ilǱ�o}��1��٘8��d�qu�ɦn̟}u	4�Ž�V�+�7�~3����١��EUѤ�"$��5嶄���$��j��+��z+.?d��QU�3!T�}���qF��P�|O}&,*��M&%����x7�@�����9����F�L�����Ǩ�@
M<�~��o�ʴ�za�PE�?�:b�3_GZZ������6�ǽ�{٩�V��V����)!H���QY��4"P0|',���+N�
�=��_��Na%��6(�
 �9ol{� �8���	��vsy�Z@d&��(#��q��&~z��^�=��]��i=�n��g?����o�O����=f9�v�*�Ԫ��� U�HNsB�5�c%��鎒��e�"�*��&B��5m9�w���XZ<�Z�,�2�#3*���p��HQugΛ�X������]���fN��q�jcX�(�{�m�ս�1���WoyX$ ����sd\�1�7���!f8iL�>�f���zR�9:
�}Í��H7�4-��Mgמ��?��M�$i9���"1���~)2&������2O����S�P=�j��U�I���G���n� ���;������L������2����P@`_���.uD6���U��]B�սT��|b$�)��J4q��;��8�
d�B%�o�������~��?���5$�i��ܬi�v9۫iG�n�V;���j����
:YOw&;�P5��Tg_�B ��v�y 뤨2:�;��G**��d]T�1�,��b�Ls��M�jဃ���+�އ�UI��`�m<���w2��n#��_f9Kp������&{�+��y�5�=��$������'���JR#m癭O�H_�Rl��^ ��`4�m��
~;S���B}4���'�y,�T�Tdڳ�q�;�ͫf��}�A�����#4�{�I.#�!�Kw'W�k��;^�2X��d�&�2���c�O1�?gb��8.Q���EɰJՋc��P���^zY�D�M̹��!8��8�P�nϐZ/�D��|Nb%m'�w���wl@�2ۂC�7��jq�k���Ūż��b��i'��pЄ�1�P5��#yT��E
�*ȵ����n ����-��b�|�n�;d�"O���#5����]-N�V�6����PWJ�(�Cˤ��<��.�5��F�PMS���L-�XGf����{{u��I�|��+�/�fQ%־��9F�j��~�<�
�u���� �t�2�s�1z��a[�o�mq��.���N!f�@��9ֺ��-��X���#�*�B�=��+.����.�览�Hbn�ߏ��;\e4}������*���0�r�B-z�AP:*5�������p)2����V7�C�ap �m�*GLy�����������)۶υ:�(<A�O$�R߳Ƿ���6�ڞ�����[A3�A�*
UHZ5a%���!�kt�:ݯlyP�]3	d�{�齕�2�koT-��;�?����Ue�N,�G�r(���矩����H�J��y�~y+[s@&�!��f^$(�ʠ���3�0 
�.]�����~JD[H�*^&M!c�_/TD�G[1Ǡ��bs�P���T0ք�s �����?F�0%m^��~rp34�jO�R��-����E�:&�('R*���~ޣ=$ѸR��C��{��܋���IWn�����Y7��^�㪅e�u�w�
"Dr��V�0�o���3k{E�G~?Ci����H���4��IN�I�%������W�C�,��Wȣ�� �l��%Cї�_Q�� t��S'OR­m�؟��� �b�iB��E��0�W1��mR��M��e�ʋോw3���6(x�;���;?G��YE��u��QU�uhr�iG�~��\��1��N���R�������֎;��y��8�&�,�ؾ~��xs�8�5R�)����ڙh����k��IoF�(��A���z+ɘGa2���Չ`"[�@��PA��UL%h���1��g}�Z��n���E��n4G ~������\e�(�{�Cp�q����j_��b���A�C�%a�?�9|(#9�l�K,�z����(z"}�,�JZV�7h�e� �9��7��[�����ҵwXj�5z�X�Ʌ)t���"~��	�JY����Wr��q��i�N\"":��و}%6��\��5�������22h����UΊǄ�֖7��yYoU��l�ʅۯK7/o�����G4�v�Ji%�82AP�P�5�Gʟ9����׫,I�(NLT��o��S��z�A
����\KBg	7� �Ӈ��C؊*�c���رjƔ9��.�ExZ����u��D�\T�z�얯{W�K� X������?�)Y���l���������]����~��_��'���G|�r��ʥS��56	\~���DC(��r�@ܱ/}v�w�e��x��)�еK~��*$b:�OX���ݚ�}z�5���]$~�ㇿ\g�~!OWJ{F�ZW(}?���[����苶�\�5�d���6�u�ǁ ��3V��@ո"�x�W�e�"�<�iΓ�S�-:7s�&���飯�ī�����˰ϛ?��"���d����.U��䡃|�24��V5aY{`O�"6�43�Qy�����5��.��((���]��h���x��8"������b����O_��+Ɇ��TI�:X9�@�kC\و�N؈��exv���]�Xg�-�@�Z��o{��~Cz>��f�Ӝ��R�CŻ�^-	���H�}����e�jh	H� �o�m�)�TI���]F���L5�1��@���Ĺ]�̞ߞc�����+��h��z�B�*"Qf��5����th@�Ry<�XCܸ�KO���!h�1'������d��Z�z�,��u(k}W:���xz�
	#N݂T}د0U(V,��1�1���]t`N2�&�JD�k3_�6h��r�"�5����S
m]Ae��&�@������KR�ֈ8�-����JO�c�-�	!���W\�_��7	���jt�R�$W�x�Z�4�8)���*4	8����_���1R�aS�\7�����L`���`��?�2�f{�P��*:Hxɠ�,��a��Bj`��%�YS��O�6so���R��cǄk��<��@�%$&��݆��	&'$����Lm����w,�  ʝ?�_�"}Jm��KV2����[���Vz�;���IHZ����D3G��Q)W�NN�M�,���+�;D�@�3��ζl	���- �aXih�H��R�m)&2H�i^`+GQ4m9�7�������K
5��ԉ�?~љf����_D"oY�lߌ�~�څg���V\x���ZC`�?��.�I8���Y�փ�i$�2 	+;�U���rx�u��}ۮ���4m��u�=.X���j�'36]��ؿ>�i��"��\Ϝˮ,�>�T�X���^�Fq,�?Bn9�7U��Mz�߰�}�n��A��7u�Q�ږ�0;0�N1
��޲<��RV��h���f%aN�?A�T��AM�����<�������%�=w{��!��峕Qh:��k4@�^���%��2��2Ϊ3֥퍘���GL-���Gq��${s���_I���1�`Y��.!�t�G����>Mf>6�uJ�Wb���&o4,�<�e����GXwI��5Mo*`�Q@ڎ�q-�L?����z��aۧm<���|﬘���J�5����*��n���ky�ܠ��)V��"��S���{~�PEܧP��8[hpX��b��bR�P#�8v�C�=#�LI�71Wb��-�+SM��p��1>e��H�m��ӱ��E5IZ�u5�t\�*�;��$E�:V�)&�o۳P�u�@Vͼ� +��`�9����*�zq�g߷��h����ƩG��Gٸ~�򚙿 �e6/�f�n�k��=�r�7�2��Hw��qL'��4CP���owaI�|�b��j>:���I�&�C��J�^����0����6s�J�o��|���i9EYJ�h;5���c05��9K֬�D)�"�m$��iF��xM��6O�b��ֱ�dO�C�?�3c�d�&VU��E�cfE��yx4_Ga�'o�?Z#/�?t�V�#����H��-ݱt<L�z���p���=��pw�lv���xנ�a�yc��_&�΃̶E�3"�������]�#���8>�(������u�a��ӫ�D*W��9�����]�ij�I�oV7*��q��x��/<�7FE� �G��e���.쬣b��єՉ��F��فl;h��6e䞼!��g�\?����%���#cE:^�O} �,�b�!����Wn&��u�.��\�#h��f���I4��~�Rd鞉Wxn�Hx���RF�l8�+�r~�EO�q�Z���43<���j�( �����t���/���N������i%S=�_�?�r���P�.��y`Z�л-���Hq��Z�2^��;9m۹�{���J��b�B,��QSoٺ��f.G-#�Y��Y�
�Liδ��0�U`ö�U���3�f�S�䘓���Nl݀iS�9@�s{�~q	o�N�/[9���n8�%6"	�s-�.�*]2��q�H�q�����Ƒ��� <���ȍR\"�@hÓ�o�F�@�'��Ը&������	��0��P4=���N���vM,13�}���N/Û�����W�[~P���k?��ˁ�ط�ȴ�����}�;�%��NJ���穀?@�x�JfCW4��VlhX�l�?��ns�Ł�M����g�r�Zƕ�-J.�b���yЎ�sU�v^^��6���ژ��}e5ԉ�1u��zp:k5���;�?E_�Jr�=�C�G��|O���=�Żd`�ZI� �jZ}ۊ~F����tr*���K{�B�xl�̵[���B_�L���p��{<Ӭy����
Ok�mJJ�%�EkuP�"[	�XI����4��2e�.�.^l'W��+)}%w���)O�j��Ѡz�>�~�m7�I������
dbX���k�Yj+��O��(6'#�nA����2>�z���N���6ȶ	m^c�*��W"��>�LnY�&T���]͚X���)�ӫX�B�a�h��ԫ�7�T;&�mӎ�����_K��~��4AW��������&l�"�?���X?}�h^H[Q+����=(z������n�&D��E������g��d��P�M���'�佘>���WvӍ1*�j��t+�dQ�]��\��'��th?�_m@��V�[����v~��!g���H���҄d�:p�K���6���Ǳ��⢴%a�u���Wܩ�d��?*-o�eEN�6j�v�@
#łƻZw��O��S���NWLPmi]�ZA��Q���p(�p���Ľ���u�K���N9�T� ʈ3E״z��п��ӢQ}>�H�"��gJ�Ls�W^�ôpv7g��`T|�u�1,k�C���ul7d7��cF����ZdV7�-����D�^�)�ʘ�_�`����Rjk���`��b�_`�(C �k�ـ���ΐ~��HW��U���S�/su�Nv2A��p�XB�S��r1�:�u�e��M�.�d,�IL�/>U����S^���8��[f���%^[?�s<��
}.�}���Bx�f���c��57�Y}��L�����>�(W��!�ݏG�0,&��f��We��B���L�Gty�L�Z��}w�a�B�|�vJ��L��T
�i�9'��6����G{�k�n²[�����#�A����htZu�Έ�N6�Z������4
!%_���"�����)����=��P�"�������m�c$��"�ϒ�n��N	�ߞH��H�P p4�� "ܸ>��'1:G!k8J�z�B\�/N�/7>B��M,nU�=��ݸ�Ѣ=m��M�ks"mA��-s�=}��Z{[�TS��_BCr�1�������W?O���pѤ˽�QL�Riu5�����r��`�/f�:��,}xU.|��@Cݕ�kw̸n�IZi�4�l���y�g�ΉQR:�EM"�@?\[Q���q���^�]��ݏ�ٜ��'�c�z���v�nڂ��%}�����
�V<�B�ų�丿 .Q�Ҕ$`�%��f�vx�M���'?��\��э�z���:�eqe��8*���iߌ�-qp�4�9��FL��-�)\�������$<��!��DԠ�ϔ�(7�͚�PVS>'�		���t���g 4�$W��,���2�e�`Ү�"��ƖmZԡ2ST�[;�4��o��"��с�.}�}�'��|�rPv�Y+��A�p�Y��;�f��B�N�B��[�Γl�kM��ݟbJ/�Z�3ڊ��O}�"b����3��}io�沮L�)�ğt�dg0`�a���@(��$:�u����g`ؑf!�f���,fھv.n�#�Fo�i���&���}$���˶*4������������<�Ȗj������W25+*.��K�jՐ��5D�K=��l(R�Y1�f=�zn�  �[�{h���ƞ
>�tA��TEh�xS�w�@�J�}�D��:����<� l�l�Fzy)܉�|j��6��Pq�_�=|�x|V ��GJ�\����	��Ҹ�+r�T�3����D��s�T��]��}2c}X�7��+E� p�6$����j���k4W>�2�n5�×�����,�/51O܋\H�"�l�  i5ؼ�)��P'�YL�M<��D����*�@��y|g�6� �ɧ��{�W�T��¼���w��Y�?L�%!n=���ES�e�>�6Dچ��H���l���Djv�+r�H�T	t�xj�>��sZ���i���e�(!a#���H�Q$Ǖ���Ķ|ǈ��J�L/�{����'���S;i�����Xh�~q��*̅��M��w��m�c>m�����*��j	<J� 4K���/��~t����w�e��-�8U��I W�D>��RL���ԓ�I&�kI�`ܣ^�^<�#5/=}��q{���,��Y�S����ΰ��6Y��f �#M�O@�'6�Hq������2�FWl@c����K90�6�^
/�EnEQ����� {}Y&D�W6�3�fC�zu��û��dbP<po�����1�g}�������x�q�����,~�x����L3�.�y���$���v��*��V���>�}�������խ;�)Q:�^�<�f�#hwu[-�Sk��E��5��"�W�_���!i� �e �4��}��G��%���2�b'$]��T�튒A=pV<Ϭ������$
��,)ojѿ��b�|�n�j��M/��ȼ��/�mrLh5�K�ϮP�jF�Wn���g��Pi�c��-��<�ܢ�`��x��6k`��K�皅K���mV�!�H�,V���|ku���}j��l9�F#�'��m�[�*Qù�Yh~������w!SlCm�W�� ��N4r'�AYm1@���k�ҒS�c����}\����1�q�W]�U����s9;@�?v�"�Ѿ~.4�Qm{�vV�'Vu�U�%R�6�9<@�ٰ�Z4�K �����`��ȧ������e��t����pN���dB��������g��[Ř���0�
Y��������0�I��m�o�Pfj�&����}B�G��\���
�-m�(o��(�K�7�	�����v~�
�c{�Ci�x-�`������S:���aӟ�"�bB�]����T��[!�"��L��A���{h�r,�r�㷠��+�Z�/��1��h-�,*����������[�S��:�i�{����y��!!>�#*��w�ov���v�DkT�IS�_ 9)�wW�"uc�i��껍����i;�u������ɣ�'
t!]������b��o�@�� <�ˠHA���[���b0KU9[���(��-;����3>����(*'_=�x���]�~^u��%��+���H�2�o��Nj��:��`]��3%6�>v#�p���,�:G���/�71�����`O����
���I*���ag�F��)�5~�5�ys�փ���Z�#�4Ԯ�
���P?HI�c�@@瀳�
9-+52K�)�+��<��{?�yH28���-�5��A��B����sF�yh��X�E���wJ�ld�8;��3��_�F�	�|_nJ�:"�~uo[ej���<>}=�>���j�+��[ f]}z�� ��+:_�]�	�'[Q͎)��x�V�.�wl�}�z#S�O�|yfb������$��[d��,*p��l���37�i�g�d��s�y�,���(������
�w@��"�4�+u��5��~��w1���d�Fx� G����)և]mw�t�6�����1����-��{6_�V�x�u[�黁��Q#���T*d�f��
\��m��3��B�֎�pY�]�|�G2���<yY38����	�D*�����S?�E�z��DW�2ԕ)S�Z���-�V�Шt&���P��c�[ԑ�0�ިҀjB�Ɛ±��0z��P�+�\�����n�O(	�V ���� p��'���9�I����0����e�̹���X��y�	C�z��mS{ u
�O���ܩ�e<ɪ@�4Ţ9V�w���
��D�X;�I��TX�1"A�UX֞q;] �R�|�Cn�P!驍�q�9���:�2X�+Z���*.��a݆?�Һ�y�<�ļ�@v
^�	c�j�U;ɹw��;6D�@�gSʵ�"$Y�}.� �(=��>C�Z��o��%�[X�i����	��,�B��yoﰁ-���MI/�ؽ�z�����W��)���Gv�7/+�/�*WI�y��{�G>N�'x�馤��2ev�z��_+�!����}Ղ�1��y��S�w`==�t�js3�;NN�Yܤ��Rg?����5��xð+���.�I�����H��K�.�9b�ʲ;��W���Cؙ��Ж:��g��9���)���`��D����o�*���́����~���_�2�*�����r��O�2r����� \����H]�?�U�3� ����\��l@�8���5V��H��ɳ��C�_� ;P��#.��S=�6�|��6�� 2D_]�dDlw�z}bt"0Nv�Gd�!XL�9�Ok����h��+r��Nh:�\~��s�t��0���Ss5���;�;�5�8u�dn5!�Ⱦg�֠��V�uE��9��y-1��Ǯ:�S��'��/xc��o{-Q��$Q>���'
N���΄���+�ǯp7l��6Ɍ�T;}� M&�v�j������4�Д������Ww�%	�$ԘXM�*<�����@:���30A�@��L�M@�
�����}X��ަpU����h�oUe���<ש-J}MXi�ȕ�v�4�+6��/���cz��M��]��������Y+�PU7�S��Uv�j�W7���@ahδ�G*���n�=���:��.��ޝ]�����e:&c:Qh �����D	�j������x�h&AO�8��p��d�rG����xV�Ffi��m���K<���:/6s_� �閑{Ӭ')��z�R%iU_��c���?���]ڌ�&����iٕt��B~�����{C
����{ Rct,��Mՙ�l����ު5�s!���d�Ua�9���2ʼ�i�n4�q����p�R��G\�I	\%�%�I"˒C���z������}vmD@v��T����B6�Y�w�"(�MU�eb@<֊���iS�7|�u�c�	+D�]�W��^�����]���E��jf��㹥'��ʘ���`�$�bM��g�����r��5�>��"\�6~+;Կ���L�?̚��b��R��w~�F���]SCا}2�t��$I�?�4������=���W�7�81CZ&�5�Y���G�hz@=�ʯ�� ��%�
�@Y�F�0�?�����|)�TbT3`MV;�# ~�Ԧ�N������r�d��@G/�;� ����A���,%Q�:����r� �^��:O��	Cs#d���c:*�oD��s;��G�<)����}�o�N�_��>2�$��	*hKL XYAS�Y#�'�@��z��7h����L8+��� ԌvTA|�iҞ5$Dr^Hy�BO�T�짇<���ז���ﻎ�o%Ķ��'�;6}�g%҉!�7q�<��W���*r�̚��C��^r�n��J�Ɇ�FWv��Tmp�s����vH��<�V	b����?���;���%����u�#T[��G�^f�]M�0���nc��c�l�g��9;���]P�#]��N���� ۟��裮�^O������G��;`�6�����wxp���ɶ�P<��d�ү����U6���U۵�b�-J&����
�8��p�ѫj0������:v�g�����OR��mCY���v	����R�|����Z�������[�Y������8���x�i�}�q7^Nl1�c��;�93�K�!`�ձM�H�f��+��]���
m�.3$oL#�a��j?�yF&U�k=ַ�'��򋲮��pw&'���򇙤Q}ȧW+��,5.���щ�V6����J��9w��6�G�Dg���e��0̸�(,;t�R��B�`
�~I��~lfs��U���t���$���""��zF�@l�,�C^@�-hљ0i C�{��1����h	��K;m�C�Ҿ�Y*SG���lXK���q���9f.ݷ\iB���s�3Ҭ��p�D���J7fu��v>&S�c��\�~ӨRM��4��l��'�n)h������}��Bu�0o�9Vy�ǣ?�ڟ�]d{�E��g��4���s���@�.V}��cy�m�����A!�v�U�SLBw��]��9JJ����4Y�0errXȠ�:(��P����u��d $�3k�϶ܯ�7��GI�,n���0�]��ߐ�HMH t܅���cYV�A��\��Q�N���?�|>;�O�HQ)} ��m�֦S!J�P�Ay���my��	^��>0@N]�
r�Ü�js�ſ��<��O��f;�Y���d�{��G2�`P�$���m�ڱ3�v𫒈�'�Dt��6<>�b�=c�����Į��q���͓̀�<#�.�)��G� 
[�
2y�Be�fx�c�Va׏����4�t|Tʞ���m�.F(�d� ��$���on֦�y�P؊�qYm��'EՍ�[_b
}�J(���� M��4�-R׷e^�K��.a����J`H��[�����H܎�PoR࿇��'$� ɆS#UD�"����_ҫ@:Tƚ4Xe�C��W�@�%g �^xW�I!�_��7r�% 5{��V`8��^+��څ�Ác�}ƃ�����x��"Om�\7s���c#�O�?���5A�X�}����*�{)�}�xoN��/6�s'eD����fd��Ӻd�Z|��G���B�U.�<H*ې�v�&����@�quڈl���>)���I���ʟ�|������:�u��D@x6���I�"t����`<��	d���Y�<o�z�F�*��4F��`�f]��|�6��tp�|��թ�]0O��}��Η�b����b�#O\���aE�ř�[+����A6�[Os��*�k�����C���U�}��	�?�k[�m�1�-�&�{�p���8�<;���ᬾ<3���G@y$A@�U��nϻ%���Tc��eO��+�5���I��L	���k���Bm��'r���\���}�L��(���>K�h���M��p���r�G��L�e2����6>u��{��ʉ�!]P��疜�%/vU�b��?p�M�c�={�ІF�XE1��q�#Q�4�uH$������8)lǧ;�V���&�f��e?J���L���t�HJ,g�m���\1R�>y��c6+KM��딎w�4�۾Ʃu9�0��@p_Du�.4�T87�cP9��n�NZ�lE���m�GJ3q��q��x���E8y���b<�Q���y���#|��/��8< �����Ɛ������ܝ��A��r���v���gZ��Ci���"5'���)vr�Og&Tl�X�a]�^6�)�	 �T��q�V�p;����)й�!�0e�)�����&�Z��m�ד���b<��������iL�5�9�� �rpv��QqB&�SqĮy���=�1{�7.>t~IX�&����%��:��,���K�ɗ�zcu~�`ׂ�K{�|gU�e-�.\�H��A&���(��Px�ZU�����m���g�f�́�{�:�0".gOO~ `8�"�MZx؊Wf�8r�;�!���!	Ht�bx<����P��e�y�7hhd5|�:<KWҊ�y�>���`a��CbVX�\�ld�`B�2[7�<���=͹��������hU"$V����>9�Nt����NEiNƟ�k�tɡ�t��b�<�,(F{Zˡ���
�ʇ��SIhs{3!/G12��ţ��)��Uw:[�8�l�+����R:������L𞂺��)]�5Q(�dR=L�Bf���p ~�s�R2|gb�[+�I�T����M�!]V8�`�����1�Q4�H��I��yI,��*j�z��ۂ�>U����x\�$���q�8�zH,#��ߦ���[>]2F��Nn~�����>nu��ف�O\�����Mء
ǂ�}r��\t�a����2U��ծZl�{�t&S,�V��9�́���ndz�;��g����")TA�b׳��?)�m���x��寃�LF<�]���z��V��>�������NE�������pʆZ�f�� 
�����[�m�Oʨ�<�j5iI�ܝ̶�q#�w��N�/c�!Y"Z���	>?M�i� c���}s�G��Lʻ&�3R��:�Y5dN��!=*cK�	�|a_��V����K%�1�O�����d�-\��p_k{��O�� A��,�s>�2��_�C׫���K��/Er~8�w���ڞ�Y�i�[ƛ^�"��:�$� >�z���:ڗ%�}��*�\!Ԇ9|G/A&��+E��޻z��ʒ"c�r����* ���/�aӎr����Mm׋�Bd�)k�Ɔ��Քy��q���Z��V����)@%&�$}�7)a���H�l���|��D�M��bt$~��d"�/Ο�4��,
뼫�E"�-�	)Fo�q��~O��新�6���������CK�1EA��3������3f觡&��ΪA\�8^�gH�ƒ�����$�`)�>�PEU��*`~>y�t0��9�Ç��׊�/�$��Y�s��cF+n^٧P^���g+e[����~���@O�DJ��J�+�C!Q�<E`P3a7Kh���q��]�L�R���F��w���|���{�/ܙQ�O3Gthz�����Tç�T?%}|�
��	�!\���(��d�2�'��b�[��TD�xF��v�Y72��t�M7J�-���"{eG*���� h'����+"p'`���;�Y�nHک+�uR�6����j��kЋe��@�[@�.Ȕ�nCt;�Np90�l5�l�ȉf�����П�J�{�oaP�|͛c�sٗ<k�f�4�<��7�>�Fmq.FW�V��d]�}z�}�$��;����DO5W��?*����`��/�'����'����&ɪ�=�%��3u4�Z�-S}�n���D�H�i�aɶ�Z�I׮XB�+s�[z��pHP��"������*�2u��^�1������*��|zx����%XSl�������8�͠^�t8��]:RN�cl��rI�8V�V[$�f�+Q1����/`� �O/��z=p��x�m��#ը��u�]m��	�2}��Ӂٍ��/:©Ō����^�Y�2X8�y�K�۝�r��RI�����I�2��J���X������9��X�vBHe�Py�SY�y�jk=�z�t��j����ic�45�T����`B�����y��)<�79$W2����|`�満C��hC~<�Ck�^.*�x閯���{���{5��M�@�mB$ϗ����H���ו;�������M�{K?\~�xAW�"!Z��wҩ��X; 
~p�5�k@'`�05���g�	�nY%?`{�l��o^��tֹQ�OJ	�u��@�>��R��C��8���N>�v�O�����k7_$#�k�F�P������;Nx���ދ�����F��Z-��ݚw��Ed� F���b��2��^�e�욽j�F��\�f4,#�$@DC��4�8��ށ���ՐT��ȑ�����%6��⻺f����E�R���F�Ꮍ�+��E��˦��Z�_M�r��;�9�Zs�{�������R�R
��S\��R���0��
.|�L��B����<Y��o��=,'9h?bIW�ã~�E^�>�/�3��N'3�D;.��)[�ET��Z����3Vb�Q�-�!�b �I���$f�0��&�6�,�e�$z����nL�h4~�T��Y�T�H0OM�y=J��,e@���nq�S��e���8-�ڌ��=_�>��k�9��	>좰�� �[4Y���N����:����[g��U\BIA�Yo0�]� f��3�k�H'��e�#uس��~W�d-�m6M������g�n�dѳ'��7L�p���+��Ðӑ�a��%��E�[y��{���w`��yCW��~�����L�/A�����"7��`�%_�Bm4|����R6�,'[ҬW��u��]�#C	��	Dz�9�S���i�1��8!:цc�U�S�w�;^~��
14�����l72GV�j�S{��I8g�!	��4[��H>�5%����p�t�R�����{Fj��B��%���T�+�z��~��[�� y� a-}B���n�YM,5�o|����)n@#���Gۓ��ē7�»a[�GdߗU2����(mc�埯��UX��)@z�M=W9�HeGȺ���%�gh����]N)]v�js�k��.�j78�IWS������LP�8�-�͏[��*���>9Z�����DC�ɲW9��l��;�Lk�X�1�D!{$r� e���v�tr��*_�7�]��,��P6iۇ#�V�sh�Qb�U�A����驆;��5�.��e
�W����|�H5�j9�e���8�sySϜ�U@���o�tv�0�`;�� Ϧi���3��z�X�r�|+���X�*�茝�r,(�w�ȳGCE6�����ˋD�a#
 �(�^cCC����Re��DE��/��?���Y��FhS�apD�nW� ��DY�Ӗ�e�I���kPk��f�M5��%Ӣ����������_�VG�3�܍p�r��G�X)�y_ca�)�iW��)�D~|�0��<�����a��?r��,{�[-���*��1��f$���������`]06a�d��v3X��$�&X���Sm�1���f\C�����aL3=r8��p� f
c"@�j�TE�B;��\�
���}	FO�e�w�1��O|�S�Q�E��I��:��I�L�ݼ@��'^p��~�����0"z�jm�K�ao�$��y�z�w� �*�\���*�����f5�� ����U���$(��B:�ܒ�iJ=	@���h��z$e��+�&,�n*�II*=ϊ@�}Wf���&le|mh�8���.�gA�r{ �`2�ؓ��O2�� �ok��W0�G~��3YD��2�8�=x�<�d�4�
�M��,@�v��af��u͆���+�5�T"���h*@ݩ-*ٛ:����z���y(�8�֓��l��LM��I�ݞ]���0�3��������t��; �^�Uٯ� ��`�ǅƯ@RD�(Z�*�$�r�H�W����c "�"���o�9i���O��
)���Sw+�;ᕷ;VO�*G�f�f�}�!wa>f�i��&U��%�����B�?n/��p���q�X6(�;�)��ʦ�ٿ�d+�C��>a�S�'���f+�A��3�!�������"��6 Q�KW��GItɂ��
�n$��f�;��&�t��f�|�1��8�!��K��O�4��7����0S�ύ��:�9e;b�����%��e�-٥�S��{�}+I��b�a��sw��
�������s�rt�/�-(�Bb
(<n�-����c
�4��j8�b+hs�P������*V�ҟmֻa�9��>\U̢�>S�����P�@z��wk2�Yg�R�6�6R������M ���l�&�e�3W���i%�i;�e���lȰ�MAO,�I��]P@g�D� d��p>�192(TG�-��繯z1.��o�j.Cr��Iq�.'tB.	w]�>���\�{�`ǋR���S�s�NՌ�w�f���U��Xc�?�5��*NalR�����"���њ�E�(�a��KW��71�oZ�8�N�0F��`���i��~�� p/Ȉ�o���t�%�;i�2���I�`��3�l�`D7q�������
 �h���H��\6S�H=}O7v6�=����0h+
É��� �Pɑehjg�Wg�P"�j�bV�l�4����&ȟm �p��):����j���7�H/+A'�b��K�Xck#|{8����V�v�f*i�c��m�۫�ɯ\��"���[Z��j�i*�Fs�d]׈�g�4J���y(
9^��L5}a��o	�'=�]l!|GI�I�v�����Ӯ"}f����-ç�LL��f���Xk;����Ԝ�=*�TK�ޱ��a�j�9��Q���Z��H��%�bk�!��5�>����%Fl�i�cޞE��{`�l�+`���x�=N��)ל�����2�s�&�n��!% ��bv{v���}� L�e[���~MŏÃ&�fB���?u�&ە�
������R��Ǿ�5�t�����Z����m��dZ ;&h;���|XH�����W�C�$�|�N~a�uM��P���,-�a<�^Tqx�{��*f�s��+q�S�л��.E󃿆^�
1��䚬e�9��U|�B�r�uJam?�A��p�>}MeŎԧp��I�מqĽQ�DS΂�!#��,������:y8X�~ϓ���0ԜB�	ˈ�#�� ^�s��Q6mZ�)����*O��2��'ӗS|�����CFψ��'��ı�h0߻1�mq>l(9&:�ga��-��+��9���J�����������Q�d�����~Ҿ�Rr����O��r����Q�Qz���`�y���=h�YƘ��=ʈ��KT�d*=o��YZM���8o{�H�W���kqx��	��t�1�~<�*�#�:F�*�D��&̲���}C�BW��$̎Q���JA�
kWU�
�ݖ�� �=6��ի� 9�P��n��n�E�eG.$Gd�n7��g��[w�B�s$�b�^�uM@K8�*�e7�{�V��l|j�R��_oy�CMlL��ǀM�8DQ�R����Ui�t,��g�0��3WGÕ::C� ��zO�t/��Ke4�	��n1�yO�k�R,��0G�]!���� �*�o/Lឳ�-���$e���ŉ��]a57�T��yA��4�Z�I�e���~O�����w�A��?/|���� �I
��"��Mi�ز�0U<�n|ƙ��S�����;�N�?�|�E3�ia:ڙb��JCK�� 3�ּ�u�K���U�uc-�%]��x }�t{���ߟd�Ó=��m��͠i;�� |�_��6K<ָb�%�{bc�������,B��&ɡױ4V޹nǖ-)S���d<�%LA��?�e�[����L�d� k�4g��e�4\��e=�)�o�H��HꚦQ�O4|����kf�i^���%�z�}�ʥ�0D�oB��t��G�mg|�`r9���~L�}��!�J�����7n ��5��F�8��]�L{G�׍'�����OǇy�x�H�"�	���{|pg�$�N\����c�#ўq�j*��=
^z[�βU��q �;��~
Z��S�򖮶G�D�8��tY+��<��Z�v3���T���rղ�0� � ��'p�U�v[�>S�,{X9P�ϯ0���L����S���ɝY�J�+H� �m�6��C�[����!�ef����[TW����}�a,B�Τ�hR��*}�3D�Q�9҅�h��T{��d�`��3�< ��:8Xi*v��/O��M���bi��p����F��>,�#��c)�ꘔ�j(볿��@����z��iYF���c:dq�̬0��*"G��\Sf\yh��k����� @Q��ڬ��]�݅�{� �s�8��J ���Z5�Sy54���Te�7�{x�>K�L�mV�]�iq�|��F�F��G�� | 2����|����=(����dҔ ��6�XZ`'��zıhdlo�+�w';��d�Ț/n51/H����s/n���TE��p������J�`(� �y����kO��}�}IL�`��ĽQĚ�`A��<'?�Di&!��$i�D��8�ygMd@tJA�D�&��'��<���U�a��%���ಔV2�H3�V�[ai���Mǘ����3�6�d�K�RC�������c�QH�>��E�>�״/ �5^�9�H�����K�b�c��v�j�pK��n��$�y1��M�]g��|�u`��钇
���F^]� ��(������x3X�J�}�iz^��5��s:�AOT�ԁ:k] �;b?�bP^��P�Tu!�<Q_�����
���}E��Z�ܧ�o�l�N��p��Z�Bl��3"�?0h���<����T�?�b�3�LbFjv�s�|���U�Ͻ�<�ս�F�����}�#Ak�P7ň�n��2���f��H7�̽k�T��J�\� 3]�*l�Q?�9!AW���q,UU��/	��j�σ=�K =ӹ�m�;e�R��cϠ�j�x��D�t�\8�r�{��y�}p4��:{�¤uK��oU}�o�2�[�M�+N>���h�%7�%mY��LQ[@	s숾�l��>�U'��H�+J�&��}h�i�|�3��>���.����۵t%��c�@c,�ϿŁ��!��&庢��5�<�߬�p_���W���.��&������]5��������?D!.�hف8��՛F��ں���5-���6H�Gh�~�,�̿qZ9�z�4}3��?n�Ok�����TZ˻a$����p��|Ah������^}W堹���!D���q'�B�����ۄv�,��8:�LD�T�苋�8bt����0����:�H���)���3i�9���+�ʗ���a;KH�J=u��Z��V��]I@��!����UG-�WZ�$Y{Tz�)��8?1D[�c,`�v[�.<�\��&��|���B�ͺB-�b���|c7�-~^X�3���Z�]k��A� ��$�¾O�hRZR�UIB^��@ZG��v�Bv3�h�*a�>;V�&W��x��m��v��:���J��@'s�U=����GD�zm1?��Ь��<��ߐ��+��v��9��1#���2�pշ���CBb��q�*����)�i�y��c�!�H'�2^]�S��D��vXpM���F�Cٻ�w��������Ě(o�j��7�d>o�}u$;��.��亮K��{�N=x$Q�ﾻ|�Ƅ�k}}��%�ȲU�&���r0	���Z"Y)7�~�GOQ9h��w7�M���/���"{w4�]g������9�1��`~�"�i h���������a�����n쇺�cCб��ˋ{�(�������Zm�/�'�t��&o?ԓC�	S��@tE)�AS;F�k�qroV}����=?�H�ʉNlH^�-��:�+���2��/��4!ӵ�ĜՐ�W�@�@��s���˾e�������v%ݢ�.%U�;3��t�{x�h����!�Eێ�;��(��0	o��_\>��*��C��hf�+f~A�$�Ktf��#ж��V��!�s�����|�0�Ōkz>{d�q�qI��\u/1�΅u˥Vm0��2�z!���>H5Y���b�z��^����S*�L��,%�E歋p-xJ�H������������d,�8j�nk�=������O�?�\��*^)ۘGF�MQ� ��
`W�Rp�2\2��K<�|��<����g"qVNb�k�"�:�P�N{_<���K�����g���"\ր[��%���<Q���
��Gl�/����0O���~z��+Y�L��=��u$P�Wy8ȼ�؃����@��x��$�9�c��9�Q��}�cn����E��]�;4۳L������Mb&��]f�uM}��\
}Z��.��E]9��)��˖�S7'���a�|P���,J(c�,�4oG�,�۞���e��6U�x/��;{SI��}�R��rB��^yOב�Ŝ^�0̉�W{J�Qzŕ�y�kѓ�b��j�4��e5��(�h�4*������.Dv"d�}�^�H���Kzq-�4n����S�)��k�j�q~����ᾱ�S�EP�qRr?z��� tE�)���)-�>*NuĪ�c�~�Z��4*���g��>��P��RD��p�?fR�6�jk�Q��9(E����=�oY�$=��f������EI����_}-�� ;�7�u����s�о���a��S�Pm����s�>W�֠��P���{?
֑���,��%��%�x֓%eMo~'m�%S��:82��F��wѩ��.)�lξ�[.�����ʵ&���IAd!ߒA�=�1�1��|H��ٮ��ɱ�њ�D�6s1f*��MC�w:Vƿ��g�cſ7nAz�/�H�Od��GRR�Ҥ��v,�-��0H�����k[���2I�"��\Ԭ�
�^�~��D����ʒ3��q�О���b���S'Z��1�$���?���)ǨN��_Q�[�=c&�#r)ڷ^lo���}�:LFݻ'K��ֱ�8�U��yKp��VEv�v�۶`T��t*�e��	��BG=i�[�A� �xu��J�-��?����Y�z�C��@O�5���m��ߴ �U�9�j���7k�)(��6}��z!�t��(x����U�)�<��	��Sh�~��1��۰�DCW��Ϙ�6`z
�7�����/��%�@oz"ݚ�(M�ւ���K[]�c�1/�n���%#Њ�] s7j��M�J F,6��]vw��aU������)��0���ɜ0𫖩4�ƇQn����P��z#73�wl�WA���1*2�E5TT���:/K��ӆ��R�x����뒿9R����u�29��Z�@�~��(��_��P��HS��#��U�9}�?��՘H�����m�lm�W���� BV�C,�i�g���b���Z�Ad��y�IC�ҧ�pvܯ��{��-U��CL���r�Q��i��RJǞ�����9y^��} �.fYSK��w�{���(�Q�5Kx���Lyu9F���kPs+H����yl��Z�+���s|�%����h>�%L ��0)����W �l�ĶS��[��<�,��:�8�
�(j(Vd)E)��}SIvPə�VZ�[��`�u��$�z%ӜG����tZ�� ��kpr|���*,����D_�B��V����F��������:��Or8J����^�1����ڷ�gj4��k0�����*u���v@a��Y-~��K���W���)�)����UG�����~0���Ϩ��C��e�eM�&ۍ�)W"Z[ѢYr4�L(�D^�Gh �\����h��\���Xv�#J�ۛt|�0���w���1ڽ9<VD#�]��MX��(����a~���q3#ߗy2�<���j�=r�27L�&Q��n-��+3��܈���&���^�d��h�K�����ܮ�6���]e����ȷ}�od(GM�Uۯ9�i���[�EeO�*����x<>���{6�K�`��m�_��,Z�̢��0���7&Y���$wCЫ�@���(�9��/�$1)_*�&y�X���;��n�~Lݮ�o�ڳA`olֺa����ڱ�]y�J.p"��&�[ռ�J�3��ς�qfCI"�	t�8�N�ڳ����h��������D�>��^�g̰.H�U:�������8�Gڛ�[�_���nRς����n�����±�m��DO}�Ў؃zk�p�{���H�9PW���SjI��`��K�U}?�&{����r����_2�!��H�}��ֽ��]��N��peIz�������6P��*�Q��V��X'{�_�TuW��P��Nk�>%����؅*�8�K��3�h��	�.6��]u��u�-��MD���7ӕ�_�E�/(%���M9K�Ua��� x#)��$g��=B�~m����1n6L��������·Փ¯0�I0Lf�DC\^�ʋ����2Q��Ǩ���X~�8��[�,��]�J��M�mG����P�����j�,'-Z�h5��8{���m�nQ���֔��k1A���m�V�X{�ԱxK�$��gݭ���Ir�Y���YT��h^ܵY��<1�o$��Cr�Q�X�x��1:&~�M���8t����8�����:��YIq~�KY�|�@�nI������۷��o����p�j.Dڠ1�4�k��%Z2�fRbo�{����A�;�߀��W��h@FԷ�0����o���[�y@p��q��.�,���͖o��r!Sya�E1~�sv"�����[�n��Eʻ:���s�@2�|Be�9�
��#��+0�0"��k���|]���yꏭfHh�ⷻ�� ���6�C�$�oZ�ݏ ���'g�%�����������AY��ni��@x�rYL�)�kZ9�i����v��Zs��BM;���1�F��霡lNx`�t���C�RZL��Eb�-)Ǎ%v�y79�W���6��ߑ#QނIv@b���t�B�7��S�2��7،�;��P�>�(�4�mSC��`������o����m�8T����~v���%1`��?�u�@Lż������rH�$�2��ВM�����g���Q��R٦��Z6�n3ɣ/��*��#���'�gX���f��.��b>h���R��v��El;�=�^,xdm�Dl��γ��d	n{LN?��(Q��~L�y)��x��~��ڥ9�tݎQD�a(oq?�=I�L�	9����@�kǒٛ��`�����e��Pg�u��ڐ(���Œ��O��팱��Y�(|"��͢뮐�;������=����+�n����1jc�p�G�� ��#�zR�{��ޙ^|�H��H8`ʭe�f˰B~�a�4d���G3�p`R�z1�NRBtR8���.6f�����w�m�/b���4�kLկ�[�K~_9����x�����~A�$Q�ga��7&����θ��ڢ~����_�j���̉�?��P��f*2߶M��U%��'���}0��-%V���e�va�^:�N�C�9���p�m�"h�(��ݭ���ѩ��A�p� ݃�D���
��x�"���*���q��.���o�{N,��e�tknO�Y�˸���b��T�Z�Ԁ��+��� ۫ЃC�ܮ:pz���S@����2����9K�����`�@[�X�Ww��^צ���P�8�Ӿ(��v;��R���=؟�����к|�_�$��+�;��S[Ci����V�1"����u�2���<����ɠ���ft�9�5_:Tb�SlX�ODc���@������P���\���!)��V�ɘ+�:����7��c^�6CE��lolim9�ՙVR|=����P�%E`��M`�YZ�.����hL�f��/�x{�`�c* 36iKm9���Ҭ1��UH�{v�t_��E�tŖm,-���
aqH��A��}{��jw�[K���I��q�:��@�z�V�ʉ�����S�5!̍r�<~0�ᛖ�u�.��$��2ׁò��f��-�0��6�9�5�F��[Y�/%4T�{ǝ.��B}�H���=�U%��B�- :�1CZ^<F�@�a�>��-���mq��Z�>:�?��Q���q�2bp�
�[G���\�%�F**y=)�9�ݕ��F��I�͇H����`� �=ѥ&'�q�\�̊7��#`������ �g�� q�3R񢬙a�v���<\p�\mr.t�Ȓ�e�J��3N����9ٔ*��\4g	Lb���2Y','I��"~�"J��8�dQ�A%��ʗv�wK&����rx��T*�ڢؙ
a���GJ�ș���8	`��C�ZEu^��ep�~;�����;[��!��'�׃9ɔ����F��]Vm[Hĕҡ{
�H��)P��b݂�`|3i"�^��*>��Y+��v��d��.d�d��D�� ^�#�&o?=e�3��8hՐန���S(��ЩT�Z�2���p
��	<��Z��B���>L���O^&U�&(ު��Ѳ�[�����Z#�5��3 ?)�L��B�X([9�N'l8_�U�z�Ca�7Y��Tjl�FG��c{��1�BbEVN��[ ��-b��X���k��m�lW�Js���9kG��cc�����ᡝ��V���N�݈x��hIi�f68�vI���z
6K���;g���^b{ɸ�d�����������$���u~0|��'��B��m1I�%Ŏ�(��!�x|��MӁ1*�h�f�M5�}�:2���잻�>�����,6�N��S��Ծ<����6̷)]]�u�m�T�a��$�Q�p�@�Ւs: Qڷ;Ps'�FY��~D��q=����_���E8Z�$@o)F t�%��s�K1
�͹+�5a~^~Z�?oӼY�
�Ԙ���+`��bm+�4��
�w�w~�.c��]D�ˀt�P����bVkv�lP��97��[�,M!�����j!g��"Oxޣ����GyMGS���>����0j�B�l�˴]�ePoO���/��<!F�
�.�W����ʥ����BB�o0�;F���
~1�}�COn�#��~ D��ѫ�E�M��b{�!��]Vfb\����|�0�	�#*�XiK�)H_�OI�F}�nH����8�(�u��TsAM��;R,�����U���Ӱ�O�2��xN�(+�vy)���=������4�3_<~n�j8�0�E�8q~2�7"+ŷ k��Y݉��ѕ�f��?3d�!��B���F:�}�/�h���,�ԥ���,�԰�i(-y�!��:]���	��C(s�T 
�M	��.~>�;�!F�.l��#u�kLz���S��H�P�3
$}.c�������M�F/���1���Jtt����z�T���K�{w��?�4³
�������$r^ͧ\�0��A�LR$��\�'TXb����u؄���I�CU��g��X��#W���4*���G��Sc�ʭ���O&�����{���LN�61ͦ���g#n��R�`��E"��p���VU���Ug䖰k̮�� � rzͨ���5��|
՟��;[h�� N8�����T�D��Fz������»{'x���_N��)8A^b3�UC�7.����u4�0䞉2s�%��B��ܷK�ذ4��l�Ts?=��ʢ]� Z|��uX�\��t�$����)Z+�3����R���m�~�-K�3Y�UӒ�~Q���fg(!7U����)uw��c���G�!�1��.dاS���i	گ|b�jt��s`�������(o
#y"�u�J#�(2Ν���>�7TB�JPW�?�VV7�wԬU_�� ��71{����t��������$�4ަP�UuȪ�e_�@��pi�IS�:,�3��p���U����T�Ƚ�<d*�����"�r��+shE��7ʪڎ���N#p9	���52 }|�7&@�z�uj���;��H/D��%A��� T�K��Co*��u�"�~^qaس�Ԅ�u�'+$�^�O+�~�+z�]��?���VKH!s]��.�+�� J�f���$O���u��e��k��ЁH���챻�'�K�[�3�i��[�?Т�~B�)���&�e<b�����>����zݮ.(}������E��+��N�«Bv��H���������W�����RÛK�C���=A�+ItA��%G6��'���j���laV+l󓫏e��Z0���4�glU1�'�~�;d�q�8f���𷍖'��޿]��:P��/D��J�fy���FS�G�vFu�=yb��9z\t�I�4i���L,�n�;�s�]}xe�F?�U���w�Mwx"?#;{�_i{�q�ٗ�_��ࢂ���z����e°���J�*��_'`V�I	�`�02�ͮ�~�4'�+��pMj�KH����+�k���
�Q;}-�RƇ���X�G�1�0PE^p��/�Y>��eЅ|�Hz��)�=���by92r�цS���M�Ã���^J�,\_�nT��Ѳv�fKr?�m��>��|#y��u�^���^��?k��i�����@#���>9$�XvM�J57�� �J��\i�lX��V�ʶ�)�ӳI�2J������5�ۗ��!��3k`��owXE��M����7PN�GZJ`�4$ۡ&�`}b���d�\�#���$[wZ�txa���?'�����T�q�ȃDA�"�>����ܯ���� 0 ŧ	��Y��]q��<�@��Q����u�溊{nzQP��n �A���̰�02�Vu�8A��Ew�"�sܫ)�Lc�A�{An���ÌD�@����_9���A��"h�t4����f�k,�L\����U�'��-��M�F��bs���	����]�}�
�#ݎ�[�X���}q!>ܼf�����aUj���Y!_�fa��i����|MS��ӫނ�A�V�խ������V�3�"��8�^"w��vS����� m���ar럑�+$�r�^u�2���0���2=s;q�������/J?�����)�R-x�4���mo�fCax�i�ڷ$���n"o#tV�h�������~0��A�X	>�&��%�W[bG��{Q�s��e����	K��xF�oR�/�[��T�M����~�+_��dMJ'�4J�'�g��8��7���gG��P����5/3�Z'�D�8/��KZJl=[b8 ɟH�5����{�9n�#N�3��X[�'�0)�v#M�����T�?GU�i��:��q �G�h����������{����Yj���SJ��}"�P�"�
W�O
�n9�����LJq��7�����9��sД�'i���Db�3j|-&�'�mA�m��%*��Gl���*��#02N�V��46X�j�k�}(j��j?IUd���.@Nʻm������#iw����q����u���k�9o��Y)��џ]�J*(�dg�/����9�f,���]����Zg��Rc�I���� EE�j���V���Pův��̥b��Q��)[�=S��,�"m����m��Q��)�&�c�,���d��0��&�ã�h2X�S��G�� (���C�M�w���ϋ�y�fkw�����y�.81���C*�+��y]I�&e�9+L2����T�B��d����o�h�J���;����3���L϶�䉁��so��~�A{i�u	�ԕ��k�[���ϝV��4�pö�[�=�JQ�`��Y�+j��b���̃!�%�$�dnr�&��!ɴ�Y	�*�1)������˩o�?[�+J5��\�#;�X�_�Q�V�#��r3G��`Ê�T�F�0��֔A�.��f�&�$���P�M~���OAa4���6׋�ڞ]��P�i��_�B�̏���`���NfǰtnS�\����Y?���GG0�e��j|%�-�[����Yz�p�u�V�I��w���$���<tr���;2���;���E�&��(����uo�|K�1r��!G$�@֞���%��3y�t?�t�О����F%�Ѻ��^��.�YwwN!-Q�ãS7�K�2��S����tSay�g����dw�h�^bX{��&��U]�3�ߙ��'~����5�=�;qzW�ţ��D���6A��&��G�B�O0�]4�$��(���W���������1��Qo�sNn�μ���5Ì��Y蹃~O�������	�F4�@ �$�Ȼ����`2��v������Wk���.��Фkv v���Ň$�DHw����R����ݩ3Y�����쀄�FF������hQ$��X��N�}���P@��n�y `f�,߀Ο&k1�+w�-�K���`�p�L\m�% Vq�5���AJie��-�<��	'h��`[�øL_,�ARKw_��%i%�	n�U�SIǑ��K��� +n �9��j�;!S9��}���P�N�_�_lw�Lf ��j���A�f��&��?M̫ba�W�!O���9M����A�I����k{�s4�ۈ��"Y�.�x�Ϛm3�����r�b��Hb/7�PQ�п�&~�Î(�����9�X�W�%1; +$��]UkNgH���%��.��8��j��Z� �������3��K��?�]I[}q�ii���_��ն%R�,���0��Z�"I9?@>�0��Z�)yN� ��l�h�d��ˮU��]�Fʌ�K0��l�b�bM�zY$*A����e�^Le�RF���N�Y�m�͆o����Ԩ/�-�e5ʭ"����L3��y�/(���U��0J�ٙ�-Sևqι�
J�\�ԋ�ubm%c�����1��H'�Ӈ����t>쁀	�f�;�iC���N�H��a/��L+2�,����zgݷa��}HY��\	�DyI}%�!>�~�ڥm�#&�;�b< :4��<�v�yx9l��#�)���b/y�������٨����d)��e��֊�1�F�y�c���*�����b-S�y׋;�<�#�a�ݠ�!���=,�����]]trJ�b�F�@Zz10��\	�|?2l�\}�y����_R��S%�5I�(�L���L�$�ӕ�#L�	
%hzz�&a��3�W��y%�D#7�v�l	����AK��K)�L}AG5'����U2۷����#�=��!d�`���T�c��X2�N?��W/z2K�ߌ��U�Pf	_�x��'\�(��g��2��f�{糇��ڮN)�e��E���ɠ�ra�7[gi�����X�	[и޺���V�A'�w#(��8y���*g�kN�b�h�f9���s"Vơ�E�C�s�i캂J�ló���ɗ���i��d�xu�.�L��CmJ�{!X�߇/�/�$P���XR�k3�;!��#9@��6֌�E�rI*��w1＄�yt�q��H�N_�[�?�_`�oS;)���j�j�r:4�������-o�� P��貹�e��p���"��mV�(W=Bj�P�8��E�y�tm�С�$2W4����~0���,C�o��=��6	�k߆�?i!�������5��Y�X��Ӻm�$/��Z+�15���6�+�L��w�&dm��]�%�Dk���F��.�w�٫���]'�3�]j@��)6x3ڤnr�w pz^D*�K�|�/
#���j�0|*u0!��1%����ŭl���P8o�Nn��)S�&���ef����m�!$���-��}CI��-;��e��3�`���E�<T2,���.N�d-�ٴ���鰺`'��$T��TUi����u�Ut�SW#n�c҃��B��x{��[~����Nt��wn�7�f,LY\B��+oe��1�
(K��?C��&N.�
��"+��6�;u�_p���4Y�h�ۉbQ���n���Q;ޫ���(V Z+�i���цDk%X*�U�li��a�}���s�I��f��R^r� �u�+]⳰)�ZKE�*Q���/���=�`P�a A�"R^T�w��1y]��d�9�;��,U�ɛ%
�%��`S�?�J�0i�-X��O(Ev�����eE��w����Y�Pg����$S�����$0���7�DbqEK��dU(���X$cf@CƲ��H��EV�[R��P�l�k���am��9������pv�ms��8Î/�� KX?�����?3W�U�촔T�3Jbb���L9�3RS��vL�J�����<Xa�$"G��$�'֦;��*Q��G!������� �޺�"l`���~�Y�Op�K3��ܙ:5l
x�Br�i& �P8�狙az�A.�*�����@L��S��=�zo!.=a�q�c�fg�N��-�YI��o��t �TwfXG��Ɣ����W��I��R֦1a[���o������jr�F��*����.��7@�Y�R��N\��qZ@�*tJ�¾&�0�u�1{�cM`y�f-��A���٦�(D�u�!J���+n�-�����C���F6�0"ƭ۳�aw���D����~��J���B^�Ռa��#�����y�������&[J�5F���k�.�h�7������lS@�#��h2��)��P$J��[m�\O+���!�X{��i#��:T��n���,��p��bj�7�Ҹ��n<�D�Os��D[�I�~(:upv}�%>��	Wo���hK*na�ƀ�!m�`�.��A�L<�d#ӡ#�!5L�L�^��kB�	��$WٶMF������
]��a�.�;s�#6��ᘚ�ҧn��f�mv�����K�����D�v:�����[���l'�\tǳ� �|uc=?����!�jϛ7=IuiЭ-����]"S.е�gf�C��nUo���q���"�,���.��Hm�H���#� mW�\��p3d�b�j�}'�/m�O�߱���g����8{��zʹ͝,d��_���x�
o�{
��Ǜ��5횲�ǋ�-rc0�ȊI���s0F��d�*�������"߸!����.���0�bI��ʼ����׈�����?]%��ـ��KP�3I�i�?zH Z����9��B*���E'�+��9�Ŀlj�h=�8�+!o=,���/Ea"�����䮈
�:rq���s��S�j��ƞ=8�u��]�)�{ �<�����IW�P�Lg<���%�cU����Q`L��v�A�oP�2M���بә�r^�ة2��IҎom?�>QUJ��{l��T�*�`Q{/�bWM��βƻ ?㞜f��z��Wa����VU�`�XvnaKae�5=kʭ�Y׀s�P�j ��s(���w��H�?R�)��i���Ί`y���f��)�'
�lE��P�&��/*�8fe
w,iZ��.X☛ވ�ڿ�R�s�HA�H�NJTH�~��2�,f�זبe��bs���n�Zb���{���������#XjI;���y�6;X���QJ�I���G��1U�\�LY��X��+���d�Ɲ���@��$�nstj��|'S���+JH.�ʴV�9+��K�mj!s�l3b^�8w��:�����4�)���% a3Ѹ�=k1�9{����eI��2tSM��/�w�E~�A=�,�� �!�9',�V"_k�ae� �U���\����	�@�������uI�BND���Cd������2�"	u,B�D����sc+�#Q.�q���E�.3���3���#D}�@�eO�4��S�q�,���'�x���0z(C�
��&���^3�r�����˽�$�>���M��񞇅���H�Y�'M��3m�Ǿ�ˮ�W �濹<L��r�֏���6����W!��b_4�$��J^�awV\M�L�a�ȿa��G�	�����yKYU�%l�4�9*�� ��1������`#Ȉ�g2��UY��C���I�RS�a��B��	d
���L�A)�u�2�s��;G0q���k-���>�o?Ĝ���9j�ue�*C;�վǗMKh{,97.���Ȩ��δ"�n�B�<���MYs\���	X�<.+қ0���<q4L4N��=���g[l_����B��xC��	��-�[��ȉ,���6�zfw�I� b`����l�D�Nkx�X��!���2���n��,�ƚԀ�eNU�Gዲ��n�p̬#��?"A�i"祲~�����
����W*�c�o�k�n'D�}g�<�42���%��>�&�{.9�*,Ý�Q��r,��`}C�DC�q�(#Bd50�.���|�:�tO���߿�&K8@-���d6�Cy����6��08:�cD=^#C���a���a�!��q!���*>�*��`1������X�E�����.R��fDL��Cl��is����$)�tu��64�W=�֛�}�9"P㌹ӍG���-I�	v�����?/a�Ԭ���6�z��1nY	f�M�Р,�Z$��-3ff>���W;;F��S��Z*DM,�`����̈�cr�)oM�D�i�O2c%{�\Gd�v���}c~s�G5u�k5�j�׃����זSz2AOd����g������[�O�x�i��Ἑ���|y��-��MP���$���A��,��9g�6*j�\/�bu���8h]����v|�x��G	q|��P���ՠf��գ��Y_s��r C%IA�	���p�Q)�e�
�/I>����gH����6��x�t���M�U,/���5�%c@R�bO����e�}�M=h�I��Z�Z�x���2��y�p�V�̠vp�i��$j7q�~(X�CL"�B0��Oe����s�
��(w�w��
t��l]���^V	���fB6���ݗ`��v��Nx_�W��&����P�B�(������٢j�a�/�#'_��=2�j*=�k����-�.�-j#�۝�eS1{	�%�f0��U=�s$����l�����,
V֩B��*�]y����ӻt��oCO���m�`J:C>�O�چ��(�.>���y���p���K����j^٣�Ľ�1<�F�8:P��,l�B���(��.�Ŭ��p~�x���I��n��K�`�B5���S�Je�C��+�#�;�� g��W�6G�Č�BԫP|�͜�jV�3�!X�Z�|�XK>�퐠b�oD�c�然r;,���������U8�.ݧ����&^�v�{)������Q<N@L9��Ƿ)R�����]�̜�eE�=۔]�ߐ� �;����HCI"Ш�pi.V�\����85�Oe0��&��<� �9��|ʦ��+�����"[�  ���JE��؟kS:i/���/�|�k�s<`���^5�X�HJ�����i�E`�DŲ\��:�i*�L��/l\�4����k�L4m	x{`6�1׾(��Ƚ�>քx�X�p(L��4$M%�����8k"�+o�{�]p:��T���C�V�>��32�{k�S��_�GI\�ܑ�5֜�)� =;��4TI�l�з��5#%��e���F�7�P5����^3R����N���4<e�aE��*��F�K�$t�fP֘�4�f:(��L_3��A�G�5��,2b�ٲ�F����$�����[�y'���|]�! ���3��0��Z�q�b�����S7~d�4e���o/)���ލ�������%���!�0�q����у�$}]
���O���<��Y2���ͤ-X��Ʉy�K��`J�����|��3��dXA�a��6�vL:ݩ@��]�C� K,�vP�j3�?�˘0�[Ť|�M�v�W+0k,���>��ʿ�M�<,C�"cN�NMF˔m���L�)�N3*C�@�2�u���>9?���2�
/�Q�W�B^���/��"ӻkP�.�@�	��`�#`�� G�hF��{}H�x���A�
GgF8Ll���bК��ã�_��?��rm5��qx �Xp$w�e�����~{4G��Q"Z��&�V��,(^ʦrw�ՀtH7S�#Y$����oZ����ڊF�2:��ڟwO���vpS�P���|�w���w�̪F�ȁ�!��Rl�B&!-��d���e��ߥ��&Kc�t۷�n�S�[W7�����ڎOc����Kym��v�t�^װ�������#
��{�H��ߍ��Ƕc���/5�Ǡ����"k������{�7�5�]�L���R���W�^�l#f��EWt��8+�k�N�� X�;��g��=�"��+�G")0����~�}�:��2(��
��*$둺�Dц����t��X��$^�<6�WNu�<K�^!������l�B�����C�i���(�`��cT������v5�$lu~���yS(����A̼G��D��R��b��s��q�F*��N*%x2�e�	ǃ+��,\Xz��Hs�V;�ٜ��R���9��v�y�;8;�+9�in������������2���`�#)����]�}��~�q�Yh��� /��(�f}�n�ALĽ�{* ��b�l�-�ᡞ�0`�+، ����b�ЎO�>�6�m;���>�Bxgb���C^���@���T��tճ�m�uƞ�[��؟�UI"ճRP2��<��(�I��Ne�5woqZ���.O�d�\��(���8��&#ϕ�`};H5�<P�O,p�n�wR�kB����N�����3��L~)���H�|���.�����d�S�z�`t�ztH�������|�yzN� Z��sG��#��1t��bIeu�ը�,����M�}��I�u�5c�dS͢�T����ަL�^�Y v��]�#`^�D$�_y,�p_M�y��юh �=X!+�ᗌ��7��]Q�������o���P(A#�r�ޓY�r�8G���RsA�e�����٥���eC9�T�_��1X�Bì��� |����̱�w8wM51���^L�4�)�i��΄���8ZG�C�	-I_��5�����'bz%�ch�Ŵ�Ə��!�m��Sj����[ D2}LRf������i!� �o��kĳ�An����6c�����A2�P�rb���A'?�KL��N����7�)�� ��j��D'LE�'����K~�;_�ץh���s6��o�ӷ0%��#��AI���/}�
TB�\e`2ʄ��yz�,���38`���ǈ�ݲ�RtX�0_��Nؘ`=�]��-V�������7�ԏ�]&E[�)9�>�y;��s�CB��BMW��͈/%:|<�`��Ǩ�ʌ���P��;;��]�%OV��Ka��$=�#�_��L�w�/����]�(��\�����K�GkF�W��0%�r���ns�)|�XcЕ�~��#d��6���J	��Ϩ���hɌ�IX��y%�(�q��~� Nƶ��,�:�̅�{�!`�F�6�Lf��Q;��H�`�v>g�"��B��B�A[!��h#^������syD]'���)��E�?ؖu�.��L:�Qw�:%��؛̩�r�n��ֆHg�3$�*�ae��jTR'�e�2�DwT	9��U�E?aÑ�4O$G��)���q�����N�v���8 �ٸ��N�0�%ٳ�I� ��g�9�u������9��aF%��X�gr����;�{<��`cf��Z��_�I��Z�%f͟�=��l������֚�� L�v:�0��u �oqr�`�خ˾��:7_�R{50g$�y)j�#�5��w�0�H3�����x�G�N�"� `���d���f�lF�,
�����O��%a�F6��3] x�N�AבW�.F�0��H�-Z��߬ݟ���*���"��qE&<�X.	�[���=ED�T�����v�=(^K����~<r��R!|����Q~t ñ�x=�Ok�o��y��~�f0� u��I�R����ÏJ�1�,p�r)��.�c�F?��2�Z����&ڦ��-A�}���%4��Ί�RηѝA�n��&Gv���I�������)���	��+�g�S�*�Ԕ��j�?��q�\n� ����!1k��l�����!��(�X�f�
��1w���ڵ�ʽj����$��2��~��\!G�e�tt-*�r�'L���9�.��;!�@����#؅��G z�2��U���duX�i��8�5�9�j�o,n�T�_�#����KMQ�Q�ViG۲���(�8l�.>0>;��n�E��<�i���PX��F�Jm5��&\���Mr�p�1�_8�0����P*>���U67��jk�ǞU��������Kx*�V�	QB��QgX�Q�%eH>7(0!�Ew���Dv9��Mni=���U�&��h��_�&ʪ��� '��'������/O�vf��t"�y�]�(�_�������s="���"~�g�O�	D#�V�׼�]Z�S�<���O��4
��r9H5��r.3	NM�#:.�+l��I�y�:e�'��"�9"8y	q?���ҋ<�q����}c�XFh�"�nG�T�M>�~*!U���v��kYPBN��N઻�Ǐ�hF����n�Iȧ����V�LHPЏMe��H���06.�w%�m���;�T���/�����@��B�ؗ��6j���w�_��(��fv�����:���Tb��^�h�w�2��/�5�F7��'X|϶��R�́���7 ����c�w�@d��Ȍݖ�1�i�Y\�M���'!�!�LY�܆d�e���i�v-�pS�t\e�Qk�[��ݥ��ܠ#$�檠� ߶8���	z3.z����Rk./�a��n{05åz��sS'�t��fV�P�¬vy�b����x���)����������/E��L -s���M=���=�+��ܮ�����}E��t�Ɲmi�X=��*`J'�EF]�-�V�}9�T�
/��M�_�Q�1�n �E�0z�:�����F�\W�M��l�3f��x��С��#�y5X�U���F���Ͻo+UanRi�6����H�5��Ea-��nA�5�h�rn��{�����j|��J��E��}l� �0��q�}�z�oS��	�X�х�^t{<��!̈���jS�g�+.��v�h	S���[��g�j#�8�Oj�+hIU�C����>]M�7v.�T��b7����5�{�jC����(䚀��#�<F������Z_sՐ0�J)�FK{�������E[
V��kﾟ5CʹB�cv�p2���h�}��,~y{���M�j��zwW_��Ł��c2cO��\�l��
]\�_}>��j�F����2�A�% ��0�@y�,���b�2hM���W���2��Ѥ;��[67]���/�f}(G"�`daU�V����?�q�����˲��C�釳f��{����<��$�:X��)ۘ�̩�A��k�[�.(�ԱD"�����y ����A�5Ϳ(�O]RGb�K� f�x�U���!��R��I]�󙪅�_�x^�ٹVI�`](L����J���z8�h#��z8�W]p�� ����Hh-rV�ޱJtkHR�k��_K&���ȏ�gS1퓔a�����2?�C����j�}d'$:��Ic��E"�Y����ԥƳ75��ǩ*&��p���m�Nh9-�wd8�w͋��E_�K]�i�{*O��3jo_��j��C9@�jleШg�6/�2ȋy��q�r	�?]�6�|�cD��S�xߔz*L����[��ޠq���z��m7����~Qv�Ti@� ��D#ݡ&>�ݖ�QV-�<8!fz�P���Mr3ᵙ�����D�ꣳ^�y�x���{'W���p�{�C�z�g�]���f/�b=����h�������fq|��C/n������t"x������-H,I��ܟ��vH�]`�d�-D@�-T�fb� 
4uD���x����MT]�a�M��2KDW5_4$�[WG�z-�[�'��bIW��Q���g��N���W���毞�R�Qk]�@��sm�}��$�]�gtL�	�Um�����Xf�/��UgwR#�C��	W#�G@ρ3�xq$B	���
$t�=ۈ��O>Z�h���a[����U+	�#cH�,��(�f���T-r���Z�0v�V[u�r �:� �>P ���õ���-�]�=�
�S`[���9p�<:r�1���S�3c�E$�
�ֶ�Z�i'j�M+��,�w��ǝ�cW������g7�w����J����^z��*�i��ݳ�x����-����T���D�[I�4~��`_��ܑ�B�I�i�\L�1�Zծ�`Nz��f�n��V�����ʱ�]a3�?k)J�l�7�,��J7�囈�A>$6j��BуC?1F쩩+�e<��Xm�Y`N'z��P-"����]�4p�ySv�P�o���|�>;�k���e��|�J��ػd�>�r|����D˷mh�PC�e�A�Z�+�����y&-�X�Aibf�1\���i�DvE�Ԁ�
��CV�J\�����N0�~Q4�B`zUy1��]^�0J`��K�a�pmP�|DF�W��1M,�z�Ė�Sɪ�N���boS��oU�� 7Xy��"�k�����.ޓ0׹HZ�$HG���K]�/zY��
]�V5���R�d���v�;�;�v.F �o���]�����Ki��/��QH�3A�i������}.^o��}�H��U��Л�Ӆ��]�����'T��N�ߴ���<NZ�g'@x)�ʧ�{��0҅aNi�ւ�m�K�5��E�4_1Z��w�H��H (ǟ�D@\F"�U7��q�4S���s���������%�W�K!�\2��,G���B�!nr�P�#��[��.y䰚{��e�0�-����� L;�i����u��"C4s�PI"��P�_w{a.[t
��A�G�.@�0��r�vmC�؂��I�������aL.��`��N��\�~�e��@��ॡ�Ġ�b9I�dL����':*֞b��M�W�/,�9n�\�K7s?99�!�����O�e�ڤ�`}����V��LƏ|pE��E��nE�bHJza9��*<߆��1�'?�3���ⶕ7�~F�T6�c/�Y
�+��}��f��R˰(Pao���|�X4]$��h
���E��z2ʖ�C����W2$'�}�N<�L�V�wj��,����/
���fj%�C,HI�F�j~�@��[���2����u��o�l�yOX��d�,�TFiB]��%��E�M��㹞��0�':�ͯ�J��&#�gPZ��}T��."�*)n'Es�6�z���j����`az��I��*X>���bͷȍ>R�^����_a�3��'���@�v�6����?,ZnC ��J��p���7K��")����ӻ��=L�G�N�N�}�.=�7�9����b؂W�L{ў\ӓ�}UF7�_�O�(y��7��`���_�vT>�(� �����H����d,|���}����k������ ��F��bv_�yk��>��꓃����S|���NesL��D��P_�0�h������AU�Eh_I�)k����z�?�:��eX��V2:R)r�����Z54�~�;��,�H;F�2�8�� L�|m,�{x�V��Y��Ğ����'��L�n�b㜘�y5����Z��@*N�����"�	���p�}"�T��� �T!�+�)�DYQ"/L���o��@�@}��T���@ƿj�4�萷5:h͙��=�����@����^A��~q�?rG�|�*GTnb���+$�G����!fu���1]Y�����x��x��;i��3>b�(���kl�����R�����U����(BS�q����eC����g\i�o���J�VA�zR����o^Y���T��[��PZ�d�����"K�*]�����b��e���K����BAv���q�<�]��O~2��AM)M���+�x�X�c<ITȆL��#�&}Ӈ%�� c$�Vx�y�U�d�G�<�@6^)?ۨ!�( {55�
+bG���8j�|��8y���U��LeiEC#v6p.��8\��%���NL*���)�S�h� �	�{�����Q��#V�.�a��^I�����jn#�T5f�Z�A4����x�hJK&A�\%�zK���ٮ�l�ٷ�PYV��9���6i"����|��]�'��t��o�u��FVs4�K��^ 	{��wq_J��T��b&���n?���+�݂-�L-���fJ9m���0��c��G &΂y,�k?�g�k���O���gw�]1&�ڞ�N:˭�c�wsI�Uo3 ~jA3вy���k�\	*�.8�j*�N7T��譚�O�/��)�i�Db���d�߉�^�cs o�]Ț��г�݁��V���*�
tv�#�`��:���<�$61�12�9�R��T�y˹�C��7�c����P�1�� A	o
���=+�E�޺V��ضӰ�q�bDp�ɞd��n�=l�g��2'�����gc�8fj4Ul��I�8r#ԇ��3�X��C �H�$�����$)�Y����t��{u��n	^�.
Ay�瀫��q ^*s(�3��X� ��K��T�`��Q>3�[GT)�<|s�se�9iʯF�Wb�]]F��o:�����u8tus�:.c�L\�`��Y��M>�T�u;g
|b�jl�$3��8�ve�W(V���U,$M\u�`�si��3�_�����f�Y���0.�����'��f��2����R�͑����i¬����h?��H�|ܴ�!�ɰU�e���Q-���M��w�w�fu�ؑr��lmŦ�<��vr0>�����	;5�:)��#��6�	�e0-�zvj!�C�m�T]k���~}��gvy)��CU�"���iXN"U����&{�BasB�I2�z�;�|��}�p���^k\���&6W�#Lm�;4
���T&'���$I�*"}d�i`�r�_�	��,na�d�Y��=f2v�ud�0U��r���'E�]�6Q���<���#�n.dH�I����<���3��"��B����B\�c�|�$������gn�ו�	���v��=�=�4��ƸWꍇ��rب���֫��r�']�;"��s➈0!��x�fO�Fd
S�M� �6�@j�q6�Bo��7�̿���z�3��Ѣ﷠���>���F/�����r!�	&�I|���Q�@��nh�P��ƞ�ʉ+L^�*����ׯѩI�++|����$�:������|���r���c�O�Ћ��y���
Q������v�V��O�F
w��;���������2��V�̥�E���p���Jlzn��#�1g`�ܢ��h=���5�J�1�O͟���[��h�"���Hێ�U���NV����
�]X�x'���mh3>������T�kOza�z� ����Q�v����6���"U3�/ڱ��k��1\���F�@M�Rm.[)�D���.;'�r�+�k>�=v|RS�`�G��(x&������3e\AQan���޾+��T4��n���z�=�}�� .�4�6����A�*� �)Z+��h�ۃܯ��m�� gR($;[���/�2����K���b��78v 0�T66��S"�@>��IN`��H�<�b�`��a��u�2��y�5_oK�h���<1m�#Y�p�����H'�`k���芰�TuR�1'�ZDN�S�y��u!7�� :���3���X?�q"q������^�N�G0\0	zw�C?�)W��{���芢�\���������?d`�����^� m=/v��F0�+�槉u��B�Y��ӔD�ʆ�r3D�-�l7�ck��k�/���K�s<L�FÕe7���M�%_n��K<;���GZ�����VQ�9��ʀ���z#�Ս"=�@!�ӷ��}L|v!v�8|@���c��]m����T�\�b� ����3 7:���&Ums�GA��dH���}��%�%��`a�PE�i�6�)źo�rgk��Jd/��	Y6�[(屢�
���t�k����cYM8�#�u�}J�����?d^�ߟ�f�P��3�������.ǉ�Tu�fc
&��X�ȡ)�ܔ����~*Xۣ���^x��7����QQ#Ef���/�6�of<\_��!�V��k���^XjY�n��+�Yr��ut�T%%G!���{|����3�2G�<Gx�O����0��XX�dP��" );�Y-�v����YNҍ�/o���V����ZՒү%+�8 /������&�ׄ>��X�nj!4;h��OⰬ�U�F��+���dU1�Β��g�VHR�X�	{��֙a��k���,E�~��V	~�,��wW���C�QTj���C1� A�(�C���t��=�����t�+Hq��r:i�HZ����</O����M�}Np�x������o�(�;uJ\AI���hQ�B�<~�|���Йl{vN�_A�R�I��f ֯��>y�(Ԟ/�d|��nZ��&�d��2h�~@�n X���M�Zuo�,�x�G_m��ҖFu2Y����u�=�׮�v�#���7�!�T6�6��R�մ9Z?��E��!M����]��\qb64>�Z�0󓤬� �OS� �.��`ԗ�i����V�V�O�t�ہ㔲[�#�~P|r{�u?�,��[
��L��<+Ŗ�LCAH����A:�H��sFO(�MN�Z�=�}[33I9]����h�����U����miP�7eG;���=P��1Yȱ7%:�im�)�يML�q�I �ě���q2t���)�J���}��p���e]��7y3��f�ͷK����m�#og�QIJ��ưv���=��O?�q�ƧDI}��Ā-ep�67lT>����lJ��h���F��l^1T�u�� Z-
�|����0����^je�u_�9uj��IeY�\��'y��|i��1���Q�'}�t�u����"K�\�$�pXo6nQ�퍈�#��9��UmШ �[G��^��u&(��#��(���u������Ţ���	DȘ�Jy�����%ֺŉ�<��I�m�������G�xH��aMS�qK(�e�E!���<a�_��Y�k�?y/�����܉!���`ެՑH�����˖�&}�i� �V��~��Q��z}���Jm��P��d��i��u �6�����7M&���j���V�|�S��ӕ8�����	�0w���P�I1�G3`8&SII���ן���4�G"C��]���W��w�u!p�m�dVӎ%
h�c|a��T�,�t�Kj�޺�2}�j
��_�1��MS(�%B"�傽�Ѻ-��^ý�-��v��(d�M�+��A�T�ot���[<��� wA̾�7)��}Ÿ떮ӊ�y����P�/1s�bq������Mq~O���E�"ִ�~t~P�d�i�ރ��Y0osto����#�,O�f,�^E�2�ʹ���Y�0#�̰Z���C�O���m�h�ΰ#iHV�-���PG�%�1rjQ�L��Y��U:�����n�³�'.�o��r_#�ª���C��h$�y�$���� �� ) ���^�3�}��lb�,N�>b���� ")d�/�WBR}�ԦF_ ޮ<N�Vi�_%��g��Q���R��jz��[��O�db�1N�L��x��I�w�%[/�d�w�{!�C��L]�qjO��d�k�'���Rn�3��ɍ��+��n4o�F�>� �`:��	G�W1�&�hC�6s��k� �QT,�aQN������y���hi����e�����*�c���q;l-�������ڑ�Ph�ߕ���#m������e��,u�����4S�`C� ȩ����l�f_�&�@�3b8*ü�pΎi��p�mq��7���$����ָ��:�Ę'�g�ɟ��i�ݮ�A䁥�s*m|�#���:���=����.�+ H�ia0��ls���%�oЩt�J|��f�7�-����f��!F~�C����������ϯ�f{�����:�]��C��F>�)��)D�KA�T�9���
����3޹){ޫ�2�_2F�:��������:PpWo�WٖߦOy[�����ʔb���b��?A��+��dY^ؐ������Z�#<��.Z}�'q�t݁b�zQ�3Ll3\�}ۆq(�@��PN}5}� :C��V��T-qP	�w	���I�9�N[�>��A�_;C���wy�H61��0����ȹ�ά���0��$E�W�Λ��@���12����1~�szN���(�y��K���:ē�2�9��}}mI� ��B�Ϣ�_ ���h�<*T�8��d��zy5b�ゆ���`���Ni���_'!����_D}^�֠�Ң�z��6�bIA�XDU�s.	2m���[_)p�z��
����P�<��@߿�/��_��~��z���^=�[[+��VoEY��JEO9^8�Ԋa@�25�Ō�:�X�H��Pi���K���j�&>��	nj�_�����ȟ�J�y�߷\��l%p������7S)�����������7��O�FP�Q�ݴ~��B���g��5��>R.	�˒��p�`�r�K��B:�y��,43���ǐ�e�'L�m<vi�O*+�e�S�����-Ml6S�`:!^��<��}����]Z`1u ׏�����e;Z�;�2���+T{����G�����£,Q���)윁`!�)]���OQ�I*6��d���ć}�2�(��ejJ�#(b�c��d���߽���d�x:x)Q���'s�\�Iφ�C���6Uۓ�+6�Np{VR��٫�Y�^=�m�����Ek
?��!�o��!��#]��Uj�+4?|��r����I�vUf�ͽ{sT~I#N���X� �/�@�Ɨ��zL��P��������ˬ�Z;oRќI��s�4��58�}:W������8�4y[�	�*���Ĕ/����H�΁��rnQO�)�,����wXu+6�T��K_�3덴4R��H��}l
Y��b�c8a�i<u�p�H=�I���6q��rV=+�}Dg�_�_k��I��P�'[r��%Bn���;C�G>�;�o���HzMzц��q�U�B)�Z7�2a-�m�Q����Cwq���ymD�"��a9���d�n���S
���h����5+��_�a��ʼ�F<b��EYOCGv��eʟ��@b�8��R�i@��X�>�������2|���V'�6�A��E�xzA��6<Nxa�EG#
4��rż'(�%�"���Y�`)���>4��:��f4\rGϛ���`�%;�==���2I�NzlSrıP��$��F�x�r����y/�i����Mw�ޗ%"���GN���iK@j�eqMwP$^X`/
���a^mi�����J㥘HW��aC�=�ɒ����Q��W$���5��U��1w�7i��X�����P0���:�2�0�eթW�G2h��V�ț~oo�P��q��X�zM)YҘ�$���	���:�%:�XO>i�w�X�8|u�]XR�T��ڍ��e������\T���3T�r�̫Pk/�n��4��s��O���:�ʴQ|�D�����c_�����4���s���L��]��V���}�y���yo�g���t�4�P�h��e�;5N�Rٮ�|VG:Dq�@�N�H�����a� e��e_W��>�v|��f���=�h: e�������v���"N����9�J�����I�]�����4��D��õ���҆lkï��Ƚӳ-�)<�A�/��E!��!�o�����]vv d���:JDV��}�V|C|���y!o�_��T�.��<����<�!
���ǙH�*[j]RM�0L�JD(��B�3	RN[	<i�ݜ˄h4��˅�M�`���Tp��炽A�K5��>��'�^����D�@Z��ԏ�����蜛j����kK��w�X���W��D^��շ��e�����Yj�V7'�h�y�g{B�����C�����2��1�����7%(���Up�/×�8wG�W������Dz%<RCj/ç[X�C�2_�?�b�`�F LL2?�l�/~]��}����;�E�%�[��{�k�iF�����
��B0�2P�p�V����֡T��\���@���Z�����5w�\���FZ�s�cĆ���eQ�e�V�4@�O�ޛ{��5Lw�Zͤ��3�-x4,Ro�?���Z�����}o����8���MQ�q����=g�ȲN�
�����T�a�s�F-1tj�9��<S�BKL`Nvg9�|%u��q[t�T^���ץ.�v����"#\7��[3�}"��O�W���u�FO��Xb]��N	O�f[<u���g��G\���	�U7$�*��|ອ��Ru|@a,o����.�	�/�g�kbh��0iߓ��l_� �
�ů���A�']&�1��8�2e��5�����,��^ꓯ��=uj"0�+��^1Z˒�̾w9`V0�õ��:J��38��x�F���+��?�JܫJcn������{s�8�ME������C0E$`�ʦ�cL�eԊb�h�.���:�w�ޥ��k��@��AH=i��@̍���XD�$��q����M!s.Hfp	��9��*�A'X�\�k�Hހx�*oY˻m۝"46�k+����Z�~�3��}W~OL�t#�~k�05{�6
Kcj���\������<���G��/<N��}��6p	�t��0��+����4�4X���i��D��:��(t�$���;���Q�f~���|#�s���`C��7���"��l�_E��<�� ����(>�� �Q#��+�8Dw���F��
�ku3uDZU�S4=�l���:!�/�b7=&V��F��FǮ�^��A���V-H��,	���% ���ch*o�t���Dk*�_�f�zw�9��pq3���Y�I ѕF���x�ṗ"u^]Ӵ�<N�Ve�q0���{���js!���i <�[�����q�o��"��1��@�!�Z��+q��q$<��?�{�6��|�8�3+v�y&/�aU��?�r��ii�"��jށ�j{C�$'xu͝�\�J���"��9О��R����lX�1ß��X�����ޫ�C��?�-I��+����Z&����ƍ� )��G�Na|�笗���*���l�����|��������=���H���\�X8'%ET~!n��D���!iT>�*'��ߜ6�=��Z7=��`0wo«�!�J��U�(Z�U<%�v��s�Pf����d��[���˯/�F?�M/j�R��?C�!N�l{3o �tO"�W����8�9eo���'�bjP)�.�A�)�Q�,�;��%�aB�y���!
hy�]6bp3;*��F��sW!�+�G�R��_ۦ������{�4��h	F�zK	�㢦��+����_2S�П�*�ѝ ��B�[�(̣%��7�҉�y"���5r(����Z�a����ȶ�B�p��Zp�r�~C�?vO�y��5N�� ]v���d{ǳPa|5]��+�i�xخ�(�̂���5�����iN�.=��fT�5DpY����ض�սl�>X%p�-���4��dM�ӹn��
��&����h���xc��ڼ:�i2�$��[����璄����U0�6�`�ӈC��=�1�ѵk���/0);O�D�/l(%3�`=p}��ĳK3�0�з��x!�[#%�Z���<j�NW#ڞ���҉#��g���Y�V���62s�cg[6���>��X;N���a���G�H��#�R꾬� ���q�v8��j��|�Y�5wu����|k�y�	:_��p +�H�pb;���w^r'��ř)�\A����`��<���k������[ƥ��*cF0`��~3[ΐ�5+dKE}~DW%�`��V�7[("�X��U*���F���*����̬�z?1"D����f2���YK=sc�_7���#�vu퓻JFQ�e�$d^(��t�θ�3GY�<z���.��WQ���i�ˌ\��͔"qygK�U�H]cm�#�zk�
B� ��{L;�C_���[��~?ms|5�)9���P�8���a��(��,�ւ� "�"�ٟǇ����$�1������$C�6���v�һ&�M�`�hh����c��k�zb�u��-]|���f��$�`~�b�)��D_d\�U�;+�~�n߷d��5�,�kA��������`IR�̋��DxHxr}(�l�VNi��(C0�p`���h ��ߍG����c�>�/�:�p���H��˘�/��vM�4��Ee��ή�Ӱ`Q�H�.I�r��hc(�̩�[rݗ�V���}D��7����:���U���Q�PVh����7�B�F����Ŷ���93�4(4½S���	�Z�2��\��G%��i�}��S����@n�٧�|�0�\���\�\�u����	�]2���f�䈮�`��W��C@J�=B��c��Z,�a|����B��֚7����=9�g\8evFVSw y��hǽ�l�M�K�!�6�.QY���b<�#��������Gȩh��)5u��+���`W��,p��K�%�N�'��w�X:a�� �D�jB����-e%w�λaQ~ýBfɬ���u��1,�t���%eCQp���R���3���v�v�l+�s(3αb܎����1 �	��+����.(ր,�uR,g*�2T��|ێ���ϭ�1R
�*���Fӆ�,ܔ4����tC�K�:��* E���L~��,��qRlzh��g��N�Zp�+Y������Sb�\OP1�ސ��*����r:�޸C`�@�n�j�>�����=�D��衭�j�SAAbb�Y#YP#�(��Q�y^j��3�i�+���P�����M�YFyXP�����g@K2}$�Q����[�9�W�&ٓ��y�]�hOQ��A����9�.�U'�������	��/3&�1�No2�K���4�'��;r/�bD2�x���t�s��&,�%We,��UǬ���H_����f�7)�Z�s0��5�r�O�.���Yu��4~k]��|�G@��nie}�ϵ�|�����/Ȋs¿˴�����a�7<C್���%0��ڕ6	�@Q���?"j����2�'�?,�ɞ���oϒ�L3s@<e�%��l���Q�y5d�ԝ`˓�����d�)��/��H���L�!��Qw��P\ �F�ErЛ�3��&P�-*�c�P{3�Շ�=���ėç����sr������4h����YhЇM�V3�����ek ��uD��/A�&�s��74�7h�G�%Q_�Mi�]	�n\��<��6
��'�Π��@S6� d@�ڗ��*u��b/���l,�~(���5�,5y}�I&:G�֢�K]8�YZ���{UV�Qhɂ6a�ӠI��w�u`���эOS��J2��
��o���[D�漪���U���n��#�~-
�,��Udk�Y�W����~2U1btĩ��a�oI3�$�_����F�����!0 n�*����lu�%�W%�c��&�ZU��5{�.l:c��ٍI��!mPJU���b[�sM)�\a������=X\U���>�����?�AR�RӐ�|�QA&T���H��x��T�Ζ�j+������(��	>H�L1(�Iӗa�~J`a�qX��p6��$�M늖�8��?ǑU�"X'�=TFp�$���9<��k����V��$��Rf�k���x�A/'e��1�A���|�r�x�cv{S4�4��_v�y�+�y��YM7p�m�E��y��,b����Z��]�ѧ�v�;D�i_�6�oKh7���#�v�%k���p��,X��z%M�:��_eX���W�,�� �^���,���yu�eT��c�m��,@�uP��|�g�Q	j*��t�:�t��Bi��٫"ڰ��p�����EP��0�~�l*��=�R�E� �ɐs[�+��66��9(�kg�nQ��A�h�����0�Y9��l\ra�����Й��Im�V��ٽ�Cm�m�7���u��N�iTi����<��Nd�/���Z��.@(�d�� ��ӽ]��LvZ�#s�7i�埻�J���A3�IJ��}2���ϻ#�}kx<�H�LH��Д� ��j���03�Đ�0�9d�
Ց�(�F�^��r��?�:�\R��+	hz+`��]z�*�>��B�1%�l[(�RlI2��w�W	���+��s�V��i�� 6��.J{Br!�)FJ�O�eg����8��J���	sX��Ey�)�6ɉ�G���b�%��8�Ywx�j+9HX�}��݀O�OJ~��A�]b�m�r`���8�yK	�O}6 �nI��b�>ͩ)����U~��A��ǂ��2[^�LG���(r'��dk���D�񭯌u��������G��a^N,p2*�",S�������cA�����'i��KFD�g�T�"���p#�1.�����,(F�]<od$4�}H]�D����J�����n*�4yh02�b��x�U���&�DJ6t��e��7V{ue�_���Ȃ�@G�wN
���'_���/�1���BU�h怑k�2$N?mr�Ƿ���0<B����EO���IF����m����IB��y��0O�LFn%2���߄eX~�4�����Y�L�����_���R�]����0�J;�bl��9��l�&����Gl�:����Tc����bt@?�m�؎�2}�}�ƻ�hh�Z��m����	c�"����`.�	�=1&�i��N�#z~[��:U��ԃ@�h���"����]w4�j_�A�̙���Y�U:��gq�T/���Ua��Hi:�-8�;�/�T��K9|��4zL
о�ha�O} �����SZ��n���삥Ң#�����瘈_�"˳�0.l�Օ!uV�լ�'����+4�X�/��]�ü��tDes#�	g�3�݊Mtݾ��D��s��%x�uC�����Ch$q��J�c���.2�4��5{��>$�Ֆ%=Ɲd��Q�6Hə�������O���{z��۾�(�vHEY|��mL�8�z�&xOL MUJ�R,k"��/��c�e��h_X�<�CƔ��_r�I�]j�G�'�8�P�"�O^.�%I��x����^� �Rf�HO����0�s	�g�
�o���2�:��&r����s]b�Nf�˶ �1�	�Mj!�9[Qc	�e�\/�z�������V�F$K���=�{ ��5�ڒ,l��G.ٳ�=$L��B_�5':��ynY������Ad\�"�;��'h�g��I>����E�_q�N3T�p���ۅ+Nj�w�)�=᲼�7��@�����%���r���5�N;S�ͥ���TGĦ��r�kx����o�?��P��נ�F�>r'ے�$NbL�n��'�ս9�	k�E0#�['�M����KA�5��	6�c�z�B:�A	��"�AN?�V͹
��/ݟO�f��=*��l�Hfq���a*<V��0����CFzhM�Y�l��,�P�/�&��.��-�Dp:�`1w�c��k��z��/0"?>}2 ^M��K����G��&��𱨠qa����K�B���s�?;��.9��F5c������uEMKx�)}�3�9�Ƞ����	1Q�KN;?����p(L�R #�v��y{���r3���FH�Ѷ�yOw��S��\-�܋�yA�܀�Ga�L�d�+8\�X�����	��ͥ���*2��Y����#nU��6��UV8��lG	�*	��L(�/:��+��KLv.�W�<��n~3�_/�T}j�8͓d�z u*M���l�T�q�u9,7�-F�Xg<4�
��	��§`���܃��
iˉE{%�#�]�t��̏·V����x�>��O�;��{�m޴�JD���:ōU��*��gp@{)�����N�����$�H��J�뢥^�g���?W��`���g��PD+���@�R�wXq�6y^�M,�Ρ��Wd�F���䳝�RP(��x�E�Ikd�o�ٹ[���}`4�Zi����~=��)s�1���U�pr~�y}�3� �)��Ǖ����Q($��_��A���uK@��*�K�b�*�wQ�O~IP�b:`����=��:^���Q՗."��_��1٪u���D��6�bW�],��c�#�/2D$o�Iz�x/H���b�H�罹��?_��@�� FP��<U�s�g�Y���D�L����~�s��"��I��b�4T	�'�!d��&6��L��e y��V�p��� ����8���d����{�c�x�W�v�N]��2�@x�ڄ�^o�Q�U�Ͷ��o�ug�Ui������D(Z� <�:���ꚛ�O�R�E���7O'�?�6YF��(h����({��
���o�*;0�ۦ�P�-"������s3�x�I�CƊ$�!pȸ�E�jq}�n�s����LK���f}qE$}ȷ?0U���F�%KИ�����}�tQ�O�D�O��� �S,Ҟ|��G�{OA�G~��ǅ2��懢�e8;��8H�d��FW���-�����ÒNs\Mo�Y܌�{��aH:������n]{��[ٔn��V�֌��J���J��a�<c:aA�Br9��줗V�����Ϯk�_(����f�U���:o�k�W���n�aLv�d���mb�טu�Y�L�I�!���'5TC>�F �n�i�J��*դ�$A���pN��@��$�*Xx�G�fL��=���6�v���%��E{ ,�7b�zB�	������9K0Px/>����\A��q�)��	�8+1�Ku�X�@L�սa�p�	�0�(r.�Ŷlӻ7Jo:�؍i���I&ra�I�C�&�!�j�īʈx��' ��`�3��AeEW��9�.�AM���Q@�����C���Y��}϶&��?]�V%�w!����c�c,-ɜ�[�̎�]���4�k81w�̌_�r��v�a�����k����*�:Z6�pe����h	]h�V�;o���-;qo��1���+��]Nz[N��ǙE��}���u���Vc�dPٞ��M��0R���zO\m��*f�oz�#ҵG�egB�;��� ��瓟�r��@���2?���),Fl����eS7A��A��9�J\���p�pw���Tb@����M ���O�?�J�1�u	����eN�lH�/�����L�������WE��L�^Z&�y��Dbdn�?����*�l�g���Ԩ�|i�ݎ��X��jգ�L��ҥO�m���c(���-��dy�K�OR�
��GK���ԥ0���w�{3��1,�|-|T��-a����4=�v�L���@OOk����y�v�����M�e���7�FU���$3�*�yS3q�o2,�J�h�GQn��§M�(j���<0g�b�ǔG7�Ec�Fy�eh�i�"_1H,�,G�I�vn��U�7	�pd�T����TlEYF`�[?�R�����4zd<m�xH�э|�#������?c�w�������oFr(:��,Fg5���@V�*�g�o�!�4��8Ky�����3�t�SS���0�D;�n���s۰�/�/�[�6����A�×�ʯ[ry���a6��oB�]o�!9Ӧ)����E�âym��(%�یA;�~�H�;�3[kL7��O|͓ �K	��څ&O��0��� Lj^ё�=�S���YHO�����0�٦$�^�����Ƒ����A2�3�*ܬ�)
���9��x�č9s�hl�ݣi���o%M�6�0&yݘ�4����T`��D��Iߞ�@gTo��Z� 5Wko�E~�co��� �	X����2�y�<V���|��� �w��H�9���J�f��~-��&��w��yk��]�����s����WqR1_~d�w�|Rq�E�"+a�|�Թ}��"�F=O�b�KT���PCi���@W�]I�mW����"�7�"9FQk���iw�"F���:I/m�K�0��"�T��zi���ܰdIϱ6Suԃ:�r�	_���Qs&��3�)�'�g�a��tew�v�i�e���j�؀S�򦳫��1�ܤ�������,!,�J}�[�t�*��:�;:�y�Q��|eE���LF1�fu���qD1i�9��.)�Z�Uy��7�BC��Hw|7���� |_��L�թ��m�����f��P�D:�/z�9���/JsRʷz�@��i�B'"���&���@�Q��*�eo��7�7�3	J��Ki���?��x��POG�=3R�[�h�YG�Kփ�؁����g�S�k�|�-�p���%j����-�S"��)�M���q0����C[K�R݁�4L��#h$�n��b:�3BgY�^<2.- 슕����:ip�ߐ�V��X<U�F�%"�F}@#�� #�R���Qg��Ju��A����u����74p��R	-�}�um+��2­���*��U�d%Fke�ꉰ�||��I5L����r�)���Q��
�"��ff4�>W2i�����Yψ&&MV�L�Jɩ�d���_?쉘���<���3�ji��+txT���0<nK7�4ҡ��R�˼�Ye��=~�6JbXG����͘�N�A���4�e%*���OYbY'�L`��'�\�[=�T�ώ��!�nT�.��)K>��|��g|�M+���+��҅
��.$TĨC��Ta<�ґ�y5�4���p�5�6Y?Ie��p��bc9�9yE$��
�� �*�@�hqY#kj�Pu���f�Z��^�xf�`�\o �[QI"�Z���PCx˵���O< XXiűG1�pgTM�0�I��Z\'"��}2c���E�!Z-�@Q�/L�h-�%�B,2䨅�lθ)Oz��"�Fi��Q���Yב]E�ƻ��������ˠ��P=TO�_�+3(��b
4���xϐ�,�+�!U�|�E[_Z �.O��h~���퐭�Q5.���v�[�|3R�n������B�� v5sX;7P�����906�{	�͚�D&ڊ[�V�O{~؈]C?I� ��a� �s�l�Rt=��_r�j#p&f�1�Gj���׼$��_�����Fƍ�ނxC�ti�-�Nx�
�rR��gT��u�$'�5Ӷ���P
+O�>;�2��������V�q~97��@~����8)C�y*3J��C���0��t�A��5i>L>���1�����4��<T�zS�,w;̞g�*���k:�8�J�v�cwt1�M'����5�?6��ٳ�'4h&{�--O��2A~���N�/O��F���1?��R��E#�F!�@䣷�Np6e�T�æK�+��̯ʝpwb��y4����Y�����-h��l�����R�
�Y�[�`GX��1`i��޸��� c��J��CێJ���yr�K]J@b�{�̽��Cy�Inn�_����>�b�����q8�o�!P����@�����R%PsV/��s|���r�(s��b�5�In�I��vE�H�q�,E"�s�Od~�ȀF�]4<x��e�+ W�:E��Ѽ���q
�	�zp�kY�EFM*��q�1�n�6<9J�R��I�W�Y{�|? 0�R�%M�a��Vc�����ܓ����P�g0ؾ��XEzb�_V��uժ��I&��ίh Y��Cx<bU�k����M��f���Biwy(y~��6NT�����}�Q��Z|���bئ^2B#T��a�,��w��B@Z0��7��8��#�l��S�� :q6i��\^��$\�z�=@�;����ht���ZL9��\�����7�m/��&'�1m�|_]oꝽ9����oP��P�=�d6����O$��������ZmZ���O��@��M�[�7Az�ֺ�N0��V_�jMzl<1R*����Fe��5!�ч�Ĉu���9).2�tug4U��$��1˭����:�q������rI��
�>4#u$������Y��ّȜ��CϤcn�n��nvy2�ָ(��|��e�r(��O�]�'ۢf]��3Z{�_9�03�|[Mh�����ͨXҶ�|�Enu��tSnXxd���������8pǢ,���pт�^>�~�c��7�K�t&*P�v����^���~dvG��֑�Z�Y(�@ñ@�鹋7��"\��0Sw�񲣣�H4Q\�b�V�I���#��τ��G:�w@���Y.���P$z��B�&E�n��|5��O���?�b�ZL���sZw��|���Up�\8�H�r�x�@� dU�	LԒs�[�̱W���-�^U�v��� �� �B��}_���AS܄�hJ*\&�K���	�~���&��KBΘ+�M�ao�^��ث,�˸�y]Gr�L���KE��~h�#=
�z�dpd8y��k�)��0Vu�b�TS�g�6H�R��xQ��o��`;L�Or�'�zZ5��hz"�19vd`�>a��&��:� Z}���r�R$g�$��J_[{�)��@u�k���%ХwY��h�>%�˯m�\�$0��7s�^Q�Cm�g�N� a��?K[+@����Ȯ|6���Ƞn���Abj��C�	i&B/?Ǖ�t[�rF���C�n�N�i,�.�S���^�yw�ݯPEw{Ū���:��!��:�n�"����m1j:��:����K�4��̕1ߏ���%a�(���V������hJ
�"����K%�nU��!$�}��baI���v`n��Q[@?�c��T,|N�өʉWt.���9�}`�t��_W�S�V|�v&كU�'�p{�-����r�H���1�[I6���rE��[%�L���1n��>l�L�[]!4F�����}+�U�C�5���Ke��w�A�{��ћF�݈��Q�D��w�z�Mp1n*7^�5�ϴ:������HN���>�`�`σ�a�\�oO�p��j6�����b7��x����Sd� ǯx8�K.��{<ҵt?�����.H��4���eA�P�az��^>j��I�X�=��{��-�xT� �����h^Cgi��B�q\)�0|�����ߚ`����*R���,@j��>��1����_��1��l&0��{:�.���%�N�f��e*r���N�:�%� �X6��X$�XR4Abeb�j��X G���3�F+��Q:q �3Ob�����M�Eb���K+ת�:*�Nt#H�8iw���>g�Bð���o}�0^j�U�Q%k欰br{��+�CMVܩ@�]��D��U���~�-�ʾ� 1:ЌS����6��	�o�/�D�;cܔ�aS�`�@�&�z�B&�C��'�g[�.X'���k����U)5>1�u�d����Li����Lx$�KM�c/X{F�+C�X�Vڰ���򽼌,րOV�ߊu��8M`9 �����3-�Ǔ[0P�t�U���!mk��$?كB�L��\٠��y���鶲�|0��R��6���	��{���j�'<8+��z	.��X+�$����},��н��,gj
E���T�aSR�BLrK���	dkl�Ƣ	���?�O���@��P׶ʟ�GMS���x���T �9��� �wޓ*��7z3�z)�̦M�GȍԢ�Fj�$Oy�	h�J���◦�Tm����Q�+�f���R�f��<vR���gbyno�2�y�w[��0�e���
0!��ɌW]����&�>#�7T���b�����dN0|mШ�_=�^Tb}Y��Rl<��dg�57�X���Ú:p���Nό���6�*9A��Z	����{�˅i�
B���cJI��/K;$�c}���.X���ъ�%�⼠���9�4�~#eo���>���]�>�5t:�ja��$ Y0�c9����r��Kr�J�7�6��#uI�w~iW�0�5nq���s9M���J��E�yu�V��Rʘ\"�k&�������b\!\��D��x�[.e���74��l�b%�
�P�xL���l4��_t: �ȣS6��4�[��d�)G�k�E̅��a�6�E�ڞe�/����5��:����2�Ƒ�!f�)K�d��$�y � ��A⤎�=)�˿s�D�8ЀASE<���a���RH\,P�s��z�|:�U��ڿ���P�*���$�[L��2x1�1Ǖ�/qp�6BZr6��d�>B�2�y<[��w܉�J(� #�X���j�c�<��D�4X���(�Aal(8��5���1[M���'�+��!�;NLq���Fǖ�2�O��>M}�Ws�raL��l	Pee`}��Ĭ]�5���\і����p��M!��~�.O� �ƾjpwY~��}s��ɏ����"(�\�Jyu	����
����d��a�["4�n��cz%�1�&�8b5���Dňk�9:`'�?��o�v� mA��hxaYۥB=������Wa�fh[0��ȟ���a�M?K�#�(&��ᑹ����\�R�U&F��^I���Ѣ[���N`�>{�E/g)c�3��`���DI��dRډ�L	h9���]����t���\�~�I���JŮ;� �&ME��ZK��r�
�vഒ�M���#��2���=�~�'N��� �[QG<���@��+�ʗ�o�{a��B�7Y}s�N}�z���T�1�:P2QM���	<\1����1�	
i�1bJ���9@��hA?S�e�TCU�?`��z�$�w����.9ξ߻��a������1Զ��rC�t�HG ?@:j��`�΁8}f��W�y��H%���Xì�zC�Z#^��DnӤ
F~�9�x�5UZ��`񂲵.�j�������L��}��WA1M�6��s���*j�2驭��i�Z���x�0ȸ^�Щ��L'+�6��6� ���hF���4��BJ�e�����=�O�q��H�
�����Z��'݊��L��@�3�����4r�?�G�v�����Q��B�":˞o(��/�S���"&
/�ܒ,�K��rŤͷ�i�f-)��i�c��z���o�����gB���N�CL��t8��Bʰ�"��^������^�p�N~K��Nf-G-:��x���U#�sl'��;�%&
@K���
�5�6�g��?38"ݩ�E2��@0��B�2�9��s?�N�8SV�Ѣ�OWj\�.T\{_���+F�虨�b�/d'a*�~\�O�\�N�ċ��Q�{-;��`�a( I5��ɢHu��|�ߪ�p#�U:͵�������h�4��,���2H�O�|�tk}B[m9=�!��G��),iD	�$���2��5��$�	��]�~cz,�|�vG�ʘ��u=X�͟f�u�)�ˀAٛ��r� c)��/ ��<\'��K&�»��3�&3WfT\M)��3�Pu�(Æ`��0A���]g�i�S��f�1]Q;ݍvc���Jk#�;�����������k\/tvz��6(-b�"�`"L"���s��y�����l7#�p��`�(���W9�������k����=��VwI��\{虍M�3�ǌCy��Z\���1�����6��H�6�Ӷ�]e6�9ZJ&E�q�-��=
��ge�a�
�#�c/�]�J���}?S����/?T�B�"�R�[+(�g/��U�� �%{!a�xԑ����S�e=�R�{��57�b�7��|?���_}=-�Ћr�Fw��
��5]b�$ҙ�]~q��﹬Eވ*��؅�ס�Pj%�hRo-kطG�΃Li�o:���fHA��$|�mK�fȻ�,�qa���RFX/}��O�aO
��8w���%�h&�c�Ki»��[����M�`t�TгF��*�#�}[ە��I2���U鄲��/nS+A� �)˗v
�����ёi ������Uܢ��92� .�����Ѱ�u[$:vj#���+�n�ڃ�0����0�&wj�%uP
��ݹ�J�Y��m���)ӂ�7]>�Gu`��g�Y�K7��>3ʷ�'��2��/����3sz��,2~�!���u9� �Dߊ
�\�">[���	��]&����a���+N ���4=�$Z�B�X]�*_\���m��B�t�����W�J���_Ȇ�oNR��~���28u�C��JL��J�c�4&���.��=�~�Qִ(���}
BȠi��0A.��J���$β0��' 6u3&�-
c��<),{��D�kY/N�x�2�PeX'���<SG��N��<fe{�U0��B2�ω��Lϵ*����4뫇�	�F]<�-k��+����آ�s���娚
փfu������nk�����w�N,j�y:���O�o��ƉTGX_�F��j�����z�&'�I���gL� b2�8�������ck�!#x��N-�6����s�5��f�t��M�`G�]�������Q_[X��Z�Bd�U�9���@����hN��#�Uu}ϩ9���ޮ`l�]-ZV�vI(WO�2/��#�����a>Z� ���z�h���\V�𹎶�7��x���y�2�K|��N���֘�;m �V�
��Uw%�E�d�������,;C��'�,T::�I'�־����8�Rɬv����i�2\a���1�N+���V[�%�Un�h�4�d��\�a���V;���y�>c�"Ȳ8K4�Q��O����b����l����~6}8沥vs/�_"r���]m���z`�z�}��
��NQ�yP�}���PZ)�-1�b�q��5d����X��[�Rp�AÅ�a��P�@Uj�u��R�L���g����x�jcj�fsV�+�%S�Ã$*Kz�f��0A�7����� "��O��d��m�FЪ%�k��kX+,������x�Hz=������8�8��Ҝ����
�����U��%;�爤�Ar�%.?���j�3��,�a��N���[�- �/eb*NVA�SSG�L&�Zx;P"�P����%>`a���.tES�zK��U�iG���=�t���Z[4RT+��1�5�2��y���vҴ@C����Űi�E$�͂���L��mμ4$N��~^�ܹM��v�V�L��r�rB$~Bc�6�G�!��y�f$���; 1=G�9۞����w��ќ�m2Ƽ%��,����ܼ�K�{�-���P������^�4� 40��g�i0n����I�\C�7B�����A����#�
\,�e|�C*�s��^L_��b[e�ћ����%ߦ1�ޥQ)� A�R�dA:<󴭥�G"�׻M��r|.)Cf����+M�J^��B>(c�J�	gS�6�l�`N�Fۿ�ɾ�=�h!�%R%Xh����/o{C�L�)F�pD�O@v���E�ŏ&<v+�&ˠ�t�"������6�s���uHz*%np ����zFO�X�
��2 /� ���T얠��P�*�6
R��M"h�x	����ʡ���Zp�JW���{��������)�4�V�N����x��w���<��p��D�7���rS��b��V������d����>����'UݼjvUo�J;_��zZ%��wfC���0��R��	���Ba��Ҁ`'��P+B};Q�an�x�:�z
�7�M�2.Xʔ��Җ�L����M�5��5F7yD��{�����c�E3.������Я���,���a�6���5K�C��:�Q��>�6��G�%?/��)9���$��Z��Ď�6��]1�;t֬$|��P��)A���� �ب����
q?�D�� ��O��n�w8�1��nB⁪	�Fj�yMn���Z��p��$��Q;��}H�2�ȁ~��6/�P3{P�UAy�J䂑��2�����1�l�������,Di�7�p�N�D�?)��;�f����P��=
β2�����W'�j�֠&���HH�J$�0B\�
&�w�7�/�	�=���1]4ݹ~ �8`D�����]��3��W����}j�9��_2����I�z�j�]��δ�,�-���0���5��$�%�9�ଠ���1��"1�h a��8�=����(�<�j���;ӱq��(�R�G��Oh�]��S2��m-)1	!o蟽�gLn��(8�t�5��
��Z��L�� ��_�s%�@�>k��I���� Ne�N���!
��.�@�E5Y���+(���m`nm�d���w���j��v��w8$�Je%���c����
}�l�s���NI �Nr����M��Ә��21��<ŏ�-f�S��s�K�=b6�ׅ(���3E0�+S}�K�<�S0�,!���?؁��l�rIOq�X��9�T�|u�V������v�pU|<PO?k� z� �s�ٟ����@p���^-p��5�ꄌG B�
ұ*L2��y�Nab4���$�2�f�V�����#��_�9��w�9HH�*�Rb	���UV%�&Ө�#yi>_�� �������XUnBS��YXX��WijA�ܗ�����K؂�z���u�a��N�B�na-�.+���Ȁ�y�}���~n��} �"5Z�4o+A�ɉ�4�ϋ$�� �K�������'���{��/��B����Z�O����o� ���YͲ�S;	o<�������q]+:9al���4T`qB���� Ϧ����s�>�G����l0CN;	���,^���48[�^�Bx�L�q���9o�}��U)�W�b�B-5�'cr��;��Pd���_v�w��T'��A�`%��+�;>�M]"�Sq&:q%�{րz@<�}���[Ҷ6~ {k7a��C���A�>pwӥz�:�Y^�5G�F��w.AMVɍh������ ��U�f��L���mhJ�P�B��X!��"%�J���Ep~����.x*�Y�t]�0��EB����һ[=��_��]�#{��'��i�E;qhx�k(eTI���.�������_��!V`��A���~>�K	Tf"'�_)S1r���$,����s="�)>�w��F~���,��j����Y�ɭ����q�(�i!yU��@��C]6vM�l�����̶�7�����0��V�'�l�=�����
���kR���s����,Fo�{��\�[�TLh�� �&�o��V�mi^�-����؊�I%�ǳ��C��*;�+sk�9Ҷ4�b�� U��L������G�BӔ��b�EAwd�\�3^�f���TM�B�7�PbA���
|&"4]6��]{ԄX*��#}��B�WD���������Q�����4��3�E����v�h�7�U��zZ��v���"����L�=�/9���j����/�Cu�~������ExuT�Ϡ��(��������g[_9�; 1|�u1���<�|	uE�o��b���JRLq�!�<&e�����N%��q���uU����-��;�e�zRA�H��{��^��φ�iN�|*##+dg�\E�ë-FDk�u��[�Kĸ`!-�׭#�}#k�Cȧ��/j�Ē��%K߮�y�� �Iה��*��A�M�����%�y\�R`���O�a�25��Оɩ�=
+��~�S��|vE�X���<m+�KKu��k���0�5߮��b����%�Λ��T�߼�v0
a����2��bG��;@�SjG�U�h2D�,[%�R�ׅE��9�4*Ɂ5E�Rw!L�IK��	�E��l��[�]�hbL���+��_u�񮽴�9a����M|V��W��7:���-Y4���^@����7���Ѻb�����t�X�}%
�����k��S<�}��5١-�5��KG�+����K��i9�o��1,l�哢У�
��J�B��k@h.�cToHAE�����OC�׾/Ȱ��'�����dZ&�q)1Q�8�������NY�9���ҒBqx)R�������ة��
=�+��B�/����j'.#�7��Σ�l�]WB"�;o��_�C;�01��iB����K�zs`��8��bc�6�D%T9^�#��E��Xõ�7�(�����Q�?b�]����ٺ�ʾr�Eg�zugi�[�,+�C��<2���	S�k1q��P�#�`���4�ՙ���^���V]
]�!#�!�oc�nHqrG�v�WޤG��Gb}=���A��^3��-�ܒ@�iә���O��ڟ"���W᛭�^��m���&��+��Wn퍕�F�ZΉ�(�RS�'9\�e�<�H_�LF"s��3L�|�0�`���fFR��w[��ʟ:�30�������ߵd��� /۾�14���.>�\�ª����>Bas���yj�����E.�p����l	�.P�X.�G��9e�|o����̛ou�ߧm=|��k�0�19�vֈ�B�>c�����s�Ǔ$T)wK�.6�E�R '����v"}#MDR(b�}�4Ϛ��8?aAZA5�x���4�)H0�ѳ�-5�a-̮s�}��$�lo<�ҝ�P�q�gM������_*����G3j|���M��j�T%���-���LۯL�͚4���djt�j,����$���艹B�k
pky`8(�'~ƍ�D� 
��_��y�[������y��+�*fnw�e��PU?c{d�*�#a���'��c'3 )|Td�"�Qp
�Q����e$�;��,r�cw>�ƲƳ�冘P�j4�˹7��e>Nf?3X\��3`�T��Еԩ�ɝ$  �����1v����8/ N~ _�-��0��x�A��1����+&��'�{�{��N�s��A�V�ƶE��\���!� ?�us-��
�M���:hQ�_������ջN@�e�	�hT�͎Ԝ�f��s
�nqx-
$8����D��B��ٺ��̉�D}A��k���xz=ÝM$Ʉ_�Ã�2W���3���5����d�5!��͐P��,��e���vLP>��EH���R=�	̜5I�@��d�r�_q���L��ݕ"��#�Ͻ>��4�nc��������k�?�)��(֏3��t��I0��!�_�3�c���sԗ��N�0�"'�	5]�Y��N�Z�F�X ��Z-����/�ev�����6d�LW�C�3�2D��Z��a�U aS�nԜ�K���n�ᱫV�I�] Ղ�߀I�$?����S�t����ں�V�ËW͜hU��#���j2 Y:o�b��:��l����m�ok���r���"�r�S5Y^h`+�O�}��{�L���h���E�(���\!��I�Fl�}�����%��[�	|P��T 9�m��EKh=و��>4,�Ҩ�P��?z.�u�h�1f�qJv��e�A��9T�_��r����T��b�}��\�։7q�1��xmZyi�*�r���x�ycF��#s�(!�iwk@���@���+ؙ�����B��Os7�-���71�}�nXF�8��) �m�6v�1��W�׹'�_����M�j�m[�ִ��j���uP�6�O^~wu
Q�ܰ���]��Ri2���ZA�㿞��t�wdo���c���� �5l4��p��FǺ0҂TO�W�賘i@�=9#�Y&2�zQTyV^��-�%�NTQL�������z��#R}�dj��"I���Ű�K�-����K�7���c�Z(PYN�|��F��������2����&U�����U��]�����Y
���UhK���]��:5�V��GY��J!�q�{j�HZv;Y�%��\�穵23�pCV�p�v��eK�ق3��rn� $�՜�R����v�4q��f�=۽գO�~?"j�T=�Cி��j�CAf~�� /T�~�o3?�� ����(6��V�Qz�������u�����|�J@k�=���c"\U��Y�r;�"M�LW�#b�3��f�w�r�f���^��b@JrMLY���y+?�W�PW}MVx���0��/�߷{�5�z��	g�9�E\��3��iV<8HQ�x��p:ך�Q���ɻ�'�%��7�rZ3ED|��P],O�*�\e��q;rk-��f�$j��ȗ��x�@}��m۰݂{��qgJ��T��F���G�B��,{�]�֌j2҃	N��C约Ӕ��B�u?����(Ѵ�BC+ ¸E4#U��&GG��	C�3�p}��id�H/(���^��~���V��^��`�m`~���L�X� �>�x�pY���\����4f���.�i�<.@ԍ�K����Wǡ6e)��} b�C�Aܮ�\�g�[ypt�^�L��2|�&�vR�ŀ.1C&�������z���<�V�m�	�tp:�
�� 1�B�
@t5�F� �?0�1�-�]zuZr�B��Tؿ��M��e6�[./��6��w���Yk�l�C�.�*���ҍ��/�뤅ȋ��ϥTͿ~�M�"*��n�wn9I[�wKG�A��@|�.wPKFC�G�<����]i2	�ƶ,�����M����Y�ʩ&�����j�`L�#��t�K7k�^D9�k,8�z*X���LB��FW�)�A�$�p���O�+�MA����5��ĞP�^|�a�J`H+��(�� �!SM�0.�z���E�y<���H��}|9n�:K���l0Ɯ�o(-ݯ�(��m<�(��RIt���	��o�w�  <�7<�:)L��X�r���Yy�G�U�����]i��<a���o�/�:N��Ya�4�*rE�W��8��G��T�[n�y�v ?B�Ĳg/�R�ݜh7,NJm����(G7he}��nhՙM��p3�k/1�@m�/��zw}���z�]M)�#�=�4�U�-Ke���\�>�x@�TQ'�V.�#/��� 
�ۗ����(��Py�ʒM����:u�K��*f��1�87�œ|%����{�x���M�fT�s��]rWk����KkK����!�DB0����"���ME���f!�J ]�8�R��W�n������� ��!ʄȡ�bX̷���>њ\3./:�;�[����
FOuI6����%�����>Jľ�_s�d*F�B ���C���b-��ѣ!��x�v�3�l�р�K ��xp�_]��H"oZ�RwӤWP�X3#���@h#�`T[zrj.oӨ+^O%�_�̓O����Ą+ �fe�WZ������g:X4�R�f��I}�h�5i��N{�M�����uv9,@�ت���eRK!$7Y#z[���(��$����/Ua��<��nvġ}
n�{���<�i�w:;�ʳe�-����HW0|�Q��ΪF{Q�6*���4���K��0< 삕-y����A��D�8�	�19������E���K��"N(�xh���|䑐4���S�Q��E�X���b�@��=�n�j�C
���Kk���i�3D��
��-����Q;����Q6���+��@OQ:5C��Fj�����?e'iTlPNtI�@=�Z�� �[2���,�M!�X�G7�:�9����b.�X���-cNV��l;��0)G�a��ɫbp�����2 �_~���31����iͨ��A�������q���A����&}t��A���|��j�B�����c�����b���S�L�����y^��7Hwl%ҁ5����}ߟ���-V h�ǰy	x���9g�"�����!TaFWBb�����=+�VkJd��xh3~��~E@��!"�ØvaOIM�;8�y�̏�;O�e�!O
YIi��ex����`1a�E��( �?�1g"U
~�;6�����2pu{�#������ H��%�_0,Y`���t�������k������^&�٥??r��ȹ7��l���8:����Kl@,��U���'}�,���+l����a�����|< b-�Z��,.��[ �)��[���g�):�1x��4x(]�0ދ�|�lIH��s�B�@>���6|����{Y�9�LrJ�/�}F��e?�gl���ٸ������I1"���jô"����D�bg�D7���>���)$P�$���YXִ��������?@x�?�T�
T�F�������r�d�Ê��h��Zp.�+�Īa�V���E���0����3#�m��̬5	��B����5���+H�(PĊ�:_!�M���%��`G7�dO��d2I��@$sC�Eӏ2����0|P���i�%�U�X"�	f����'V��-�!Ț�R�\��@�k����R�2nђ�z�P9'~����ud[������-�Ў.�Ð����q=�Y���%����q	�� ��/=�6}���	M2p�^1p$y;�Tz�,Y�ӓ��r����T0��x��Y��%s�/5��08�	��J� ��֢ �ݡ�]���(��(�!L���qj���OOY��m8W��v�0ج@������Ђ����������i����~�MG��� Gn���&�Z�0Z8�X3WW_ݧV�;I�1��>g���>�/��#���Jk���μ���RCn�l��ۻ=ć�Vt]B�]���ǖ����.����^�X�F�z�䮫N��C���T>�u�y�GQP�FY��v�q�oɞ�!�z�f�]�ݨ�Ӱ�B��Ң����['@�P�ǣK;��6	pjfmN�|�J�{�J�"��4*bhQ��.�M�z�e��j�M^��/8O$`bu6�%N����Ex ��3�	0 f�K3��vH�/|�D�"������[x��	O�4/��5��"��P��A`ٍ�c8��-\�e�M�&w��� ��i�Xd4u^x�[�;�ُ������t7��+}cQYSL�t�*M`��G:�y���rH�E�1rcE�w����6/F���=�4Q��4"o �}��m?��Z�hR�7��L���H���:Q�haJ����o��'Z��K�ʿ��%��x�`���d~`��@����B0&��ߙ�V8ڻ@��G"�}kA��!<TB�_E�Z66��	��#�urą��GCDw���,�0���E!�
+����^��'��#8�Q���g���b;)s_���=�U��X&( g�{n��)�D�a�Z_�T�3� �岰|�Rnkv��p������׌�Ge}�E�C�O��7��)��E^�\��2�(�EMPw�^�D����W?{��E�k�� �@�Q�J�
L��^�t�����E"�LH�����o�X�~7�B] WkuȲ�����H�%2�=��A!�̠�����Vn�Q��,�^��'(�?�pquB4Q%tˉ�~L�T�V���Q�}_�v��c�TY�V�[��L��H��W"ƐN4���F���e��K6�[��Ti�P�#`�{�"�vsI��Q���{å��ʗS��e6��ଦwV�-:>y�"o5S?�Ev�Y<-G$xb����|v�QͮC���I�N�*�l�Sj�J��A=��s/��; .�s�D�p� lJd���D��0��|hl��w&he=X�ۋ�{�vP�-e���׾����N�P�z|T��-��}���=�NFW�?{�1e�A�i:F�y;�gL��ǭ�w&2���k�ֺ=��.�X�y�4{�YG²��0.,Ooo�������e����R������w��d��_����ry��z�w �sy��o�t�P���ֈ�4���Yl�m�s*��c�*L��aM7W���<ƫ���^K����X٦;����\m�o�H�sB��~��]~�|��!��}��?��g2�7��]�"
c�|G3{�\�����х��h�H�!�ڕ�@� GlΦ/�fn�E�B����::ꈽd?��A�����-��(����#��r�:ش���?���E+2�DxP`%(�e�q0�X�5P)�2/��`xH.��VHя�����=;z+"r���jp�d;ܹ�ei�֊�LC���H脚Sz�pi	$��`i��x��?D��H��=�_������j�(w��4��"��� ��h��Y\l��z˪2�_�����"k8L���Y"ќmm�>���[�)@5��>����z�� bZu�ؠH�����F��⠰a8��b��T�����Q
���r�8�S�s�]���8���?�`�;N 4�7l/U]}26��V��/f��RL��)����?ˏ;b�D5����=��Q���.t~�ޚ΢�J�Z���o�����B�*s�^����B����;L{���#��g�ūf��r荒��bև��7Ȋ�4�Ė���~ޫ'RE�֤=d�mؙ������r��Sy��NW���`1�$8��/}� >��٭�����J�wW��F��ڙU.�����vN:����9��BG�y�Ʋ�G!�*�ӟL'^[�l�k����iNm���d���Rte��D���T�H>�f=t�j����a���R}+Zg����t�sM'���;��[wf8���$Д[��q��N-p5=�E��đk]�F�m��on�&pDV�}�G�D��,���'�K�
���98�.K���b�5�3�P��<6$�5��z�)8S붌��HX§[�W�%���\�&�oR-+xǃ+�g#P��j�$�9�J�|3�����n��Sx0/RN9p��\,Z1�������X��X��mg-�k���@�X���xU3{�o_���]�了�}5w�qi�t�6}8~�����s
cLo����qj����hyn˜���ݚ�P�[�`VdM������`���e�V~,�C=��pzΖخ�h�72̛cߎ��ŧ�f��Z��	�	^���P�쩾��U�|��r�[��T-:rC\ɇ�п�UK�\��-��O����u_B�rEy�5�jx.D����^�M�QM�f�)���xSG[H��aiQ��\�2�O��=�4��	1��#9����1�M��]��[�g>���q^������'>R��ob
��g5k�#�q]ڛY�"^�$���#|�EW	������8%�3��;��]�B����aX@'��*"�m���,_���/|pFO{8�-��XZ�F��=��E��Ni��g��6TD���zavn�T�>k4姚'�D�ͮ�r��=L���zR�C�R���z����s"�=�aW�����C��~����;S��pJ�_����;˩9�4������ 3�6=�#wt$wC���t�����ò� ��-�s��d���#i�$�d�3`@�������������,N�aR�K�4�e%���q����0���ۡ�)���
`���
�jJ�Cs�L�+'éJ���m�e������@�aZ)��"�}���CћYĝ8{L�Cq�ݎ�`߭tC��4��y�� ���	ވ����Pb�^+R.��0̻��i_��,/�P�r؞e���>]_9RO�tB���M�;���נ%.����%�췪M�K[z]Z_�Ѝ��]�	v�!d�}�� 97�w�K')y�31��ԕ�Wj��}a!���L~:'�S��)5��a�Gi�/mC�v���}<>9{�O](HʭaR.Ht %L`�?��5k+��_"u%��^=������g��N)0,��b���	R��/��-����R�(V��|���-�y��~���%:_�����0��+����ŋ E� x鲎N��t˔Ë���}�uv�#���? �V����ņ���M�����X�9S��p�4��g*R����3�����^�n�����v�����g�\�W��^?Uk;Ԫ/~���1Wh��!B?��q���E|fn�u��C�\xe���Y�(�vy+�5s*"|��S7��"�%���	A]&ڼ�C���.u��³D�~q��Ki�)����
o)l4z�S��=W�s/��1��Աd��Y�?^���+���2te${�X ��ȃ���8���'rDڝ�b�䳉���h�N���Ždz¸{q�^�m�����)�^gv�"#Ee��4�\t:���D����D]���4�D�;�h*v��;ǈݯ&��{&�6w��C�l��Ӆ�����B�A�M0ۃe?[�ױ�ߟ��򘨨���n�f �� hq�i��Yև�C�)ڶt;7�
t"�	w.
q�Rj��T�"m5Ǻ�t��a-��J��{؅o�O��:�V�C��F�cm�5���*}SSh�A�c�k���+I��u0Ca�����OK���0�厝�C�Vz���Ⱦ���s��1�%��ԥ/`!�$٤�k�nqmL��J�:�
>6�˵7�@��3K%�:��C��[H� A��4CU]��Z�Eod&��4��,i7��u�M�dpk�o17km�R�yq?S�Sn��[+��v���\=��`qYZ����j{�gB� M���M���n� aO�<t�
VI��y �h&nj�4tA�>�}��h^P�z�/�V���F�:�����j@�Խ�wy5�:���I�V�3*F���^b�F;-�Ə3p�m��TeQ=�.��MU,��PO��P�k54��d,��>u^��?u�R�\U�B49�zW��a�^��m��a@�,�O�!Q���� KT��{��&_� ��u!˚�r�( 8 H��4!�Y���"��U�n`���7�!��dhܢ��LRx����ck'�wz��c�͖���;������2���J�)�"h�B(c�4Ɂ��bA�%t0W�0�ii��H:��pn�so~ƀöz~]�x��ŌF����7s��>���)����EY��Dl� g]>�\�0Ə�sW�	����ް+� �r|��g�Ȁ	N#� Q�:��I..�e�_�����R��*�
�N�������2�ƿ��h+����l`r.w��M0�;�FE��#�w�Q��}����+ݳ7eo�,��0��:��eXk�Y�ZÊ�]�S�4J�y�����+�b �� 0]��l��^�,�=(%Px��G4MC��n�i�򁯵������n���I͊�	�@~j{"q�^c�g�x����r  P?L�Z�:2YŸ^�|�G�4�r�a�[��6����N���9���z�X�ĭݨz���p�o��NQ[0%ĝb���gm,���b��:��*b��p���(��^KV�FV�����$\����{mU�����7�녹F�Ff�g�T�Y�2fDX#���=Xe�a�Cb��ؘ0�z���8 �*Mb� w�����A1
�`+ߪ�_C���_O��4�ۢ���:T	uY$q@�b8�ٛd�����J�~A��ov�d�*Z�(�U� ������.弁jQ�p�aI"B��*�c���V c�~R���3�fX��_ƃ"�"�f��:~F��[qY^�<!g�jccy,/	�µw�ݟ�S��J���;�(��2��cM>����g{�d'��ٽv���@i�7�Z���R���w��S��и�y�⤧P�5¤h�v0Ǳf���j�3K~R�i�£����4̈FtQϫ1k8%� �jy�1sʓ�˹t�ľ<�wk�� 4U�a�Er��T�q�e�-,I��칉�2�p}%K��޷�����mM�r�U��r�w+S,�序�������PTCt���o\h=;�<�Τm�ǻD���Lĺ���32��r������o�57)��˰�.J�/��MU�<�x_��$�hD���4���v�VBcv`! �4�VJY��s��'�l�H�c̭su��Ӱ�*�|Ӑ�E�sNZ��d�� t0����+���M;��S���lk��NaP��f�އ/5���
BDߛ�a@������}f�o\�М����mگ/�}��@󏗌E��
�P�S�f�v�{��ጮ��Бx�8F�;W���b�B��^y�+`��c'on�<����:S8����z-F��W�"�vrȌ�������y����͒�%j9���e�&�@2V�	��ޡ����Խ�sٮN�>�����x��*/D�ɓ������f�в�v*���_E������3��k��YM$�{4�"���]ԅTC�,���!���5H�B8s�����������U��P�K:��&��O�Pd
׫�0�!�t��:�徱�\?O�������I���y;���N�ןr�?����Ρv����"@���Sz�1̄������"���3H �M�)iG�k�x������R��zC��xmt?ز8jŧ�j�����K�hzm��R��N���b�؅rD&PM��l��kv5*��9 =�	ʓ\.�xUo*��}�eA���jiԋX�����9�BLI#4�\������k<�j5�H*]V!eR���[��$Wg-œ�����9@� f����g�+$���R�<�|�g�u��� �9��M�q]�q��B�\�LY v	�A����m����p鋃�`��)�=f��X��e��۷ģR _
f"�L>�ʰm,@�v���Nʈ�2���j�dω�Ȝ2^oJn��1�j����=���A��e�H4���%��@&�a e�I�� @�X�$���o��@W�`�h��}�p�zW��J�hVp��{okp�U>-��Cɍ�SYe���/V]�7vL=��x�kAb���ӁΙ��	m���f��@��j�H�]m�v*
P�4�`_����߸���$h����k�$�/����i:0���P:���l�C12}(QIl����pg�� Q[ǜqϩo�RL���*PF�\��\��E	u����n��3(#Ę���~��k��x����0�=�y����)�[|��A�o�hRzV� ����-�eW�)�4�uD{�տQ�}ٶF���� �=5�_ �y�����'��O�uX�t�R�c:4,_���n^����Y�gP EB� 0�D�I��Y�B�A4��mۗ�v�� �߅��O0�M�vƝ��2��]�+&�����;�Y$�Υ(4���P�����|X�M���^�3�(��x��*�MG?�fю�Yh����ޭ��(V�2�����
��;���F�1��ӯP$�"�6�~Yz��XS���x8h/x�6�OC��+�<����k��%��L�]dD4�&|W��a"$�9L[S���g�\�~���m��ֺ���K��տ^WT~"t���	�yJ�$^xV=�R�4W�<�5a� �8�Wg���6����T�b��^7ݪMvd�"��!�L˭�W���P ��D̅7M�rRaA�bKȾe�KLH=��x�	������teX�*g��.H�d�i����T�}�T#E�G�Z�ƫ.�O	l��N8ߔ�h���q^��x�p�k�wb<���g�6Aȿ{#s���w�:qN�U�ڇ��T�@Po����8��_##�X	��s̮���W�h��}(�3�2��io�F�`�w3��P���Λ�>7��"���hn6�K���h�J�e6���u�Q�svG��60[�B�o�(�/��ui:�#ȷ��_P"w�>H�v/�tT���̲��J�DxQ�0�!0V�l�t�%�{q�u!����zP?�<}�Q@Y2	7�"ε�J�e���.�D�8$�?��>*l�Q~��Ű�����I��Q��vv�WT�dcǎw��I^���4/V�R�Ʃ�I�����-�S@n��`3����r=.JDkPuB˰m_F/H;9�iMGqm*���0�MP���R��d�DՄh�p�������c���ŷ����D���U���}4���H��F���R/�J��%�\2;�
/��{H��޲�4C�o�-᥃�i�F�J<p��|�B�CW��9o����Eу^U0�o�L#��~DlS`6vq�9�ځLƨ��,���Rŗ�CC�=�K��x�Q���A��B��}�be"9�����l������
��Z�Aw�}l�U��..\�[���]��{�M�a��[�Y�S�5k���ύ�RE<A��B��V0lIh���dRf����c��e�z�ֹ�ҴEkdljqOK�
lnEi��
.�b������Jo����~�2˺�f߱T��p���ۇ�����\�ޓ�T���1�u����&�U��;r��<O�2�h���
��3�(�s#*�z���W�?�L�#�OjhzDs�8e�G7�6Y��0v�n?p�~m��=�1+\����f9� s0���+�>����:>W٠(&]��"�MK�ch��t��vD9K�0��e��j3_��ؘ�{k���0U��7a��Z��g��k�&�ī���}���-�#�}��AF���� v	�?�,�X�j�����5Y��'��y�8���y�|�~�|�:���~Ʈ��lj�L��%� �wX�d��w��|
�p�Ma�0�����VgT{fm�9��[�Y-��9���v�m��ݣ�og>�ܼw��R#�o��q�ȫ�������Jy ��I3[�V���1�;6�J%7�f�^��8�(V�7�+9������UW��c ;-���B��-^�z��@|���ۄ��H��*���%�P�n8B&�:�F4��2Y�y�2�F��5h��S7*�6d�S����aſvg)���6�lj4�nԮS 	6��S�)�,�XZY]"f�/-7~��j�KөO�H87�
ѩ7�ڏ�Ǆ i^��92��*�Ƈ��R�eo����_��_d��.�)/��J��"7���N#kJ[�r=�q��s�q/��� e��p >�µM�#@?=���H3��^�
���bR~��ש�PE�����ϐ�Bv��b:&-0��/�s��E�
�� �+ٯ�/��r��7j|/������1��E��L�Q�vnl$%�/a���G�e���v8�vg|�MI�\U����-`�r_R���]阣tʔ+�	��L�����ƨ����N鹧v�Bo�d"��F�v�1��P��`��l��
V���O�<#ڲ+5��y*�e_�@'?��2F�l%d�a8��e����$�$Å�',0"�m������`CJ���1�1ֿ��'�}��Ƴ��aț�6���Z��Y
�^�=& ��<Z4ݟCP�i6]�<�)a���7�|�<�r�� ��`6<)�}����x:��5E`����boϞ��.p�H�*��<(	P97�%5/����)��n�B��`��K٧�z��֒�A��6ۿy�:����b�#T�x��]�Vj����5��%0˥[@N�	��>�D:A��g�^Sˍ�Q���Eċ��Ҹп~}�DU$\+�F�/ ��V�|�6�bV iB��/i,a2�
<!hvP#�Z��Pߩ��d!9�1�
/�̥��k�G_9� 7"g;Z��n6R88��;KYԶ��5Ɏ]b�H�za�����S�3�!��*+L�EIr%�O�4�����E@\�zK(P������P�Tm?�yZ5�I/�o*���d��y{h�V]_R��R�[������3O3B����L̗���M�Vi���1�#Uq��?
M�XM8���"& =������g{������N�^-��<�9<Y�������9bf�E�Rcѿ �yA��!�@�nؼ�eЅʫ=�NO�s K��8�xրMȗ�XV��f@5��+,�f|p��=�
���t�ggT6|�_i���{��W�z9���#�~���f$�FMf�/ɮ�Qd���{cA[���J��B�iÎ}V2;�rMZ���Y*h-0J���$1���`t|�ƣ�'k�&����ݑ�vM�k��c`}��HYH�L�����C���8zo����\�fN}��x��$�
���j��C j�D��6gB�����ӝʜM��@߅�r�QD�O� ��c�O89[@�ۋ�:h���)�*��qi��y�Y����$/#D =	ʆ̳�5������
u�I��V�E!��� �4}�tM�g���X�Xk���(|�)����F0���D��S��_�	g)k�+N}�9���{���^�j���V�9�F�m���@S����?������1�j�9��nC�B�d
����-B�\-VP�h��~ C�U�b[��'\�L�0�뉿�kr(Wf��&y�4�����Ra���푆t����S����8H����)����x}�t��kU9���*�����r�����G���:<n��sۆ:�k�Q����"��E^"�h0��(){^1H�=.�0�("�Ԏ P�gJ)v�׮�^u��ߛ�t�Ψ��]L���\B[�k2�:L�� �)0����P"##J�t�aq ����/z���Xhu0�"�S��w)���������#o�9b�:
W�x�dt��O��x��:�w� �O�����x{��d"��tAp�/��Z�j��k�;�HLw6Dr�-�r{x��Ůfƣ�'r�D)0G/��G�k��Py#��*326�<��'��/�eF��N`� ���u�﹌ۤ��D_�L2Sl#����T��Vi"��l����@���H3y"���3r>G^�7����m��v|�;`8ˊ�r�� 5&6yP������`�����[��i�� ca��\qNt�;X�U����=&��-�A\)���[�3�)���[c2�Љ���.�c��VD��e���a2�mir9�T�.��Id��c��)~��|d3�u��; �9�����r��]�+tR�G7�Rc�;�oN�)�R��K�!q��W��� 9���t���)����ø� k�l�ǖ��������&����%p��櫋^�0�不����}| $#ά㐩"��eK�ں����%9o�Y�+�I,�M�"�?�\���_g��w�0"`l{�vO�����YY�A�4� �8wf���u�{�/%���]kԫX��ۧ��Ͼ�g$ чW������9Dv:?M�x���4	�b^�Tݜ�"E�N/�2��/�.��ehC�����D0������P��3f�����9�����C3��>5�Z4�K�8��D�4�z�GO�����e���B8)��v?)�����YnrW^+�܍e����P�-�Տ,p
�������iرa��Ϻ�@c�
��N�ܩ#�����;�μUx���ȊZ���ï�E�h���?[�{�v�G�N�@�.{��B�x Rb[������_��-Y���}���8 	>54�wA��[5{�g�D�>�3>��+/�g��j�lҹZJ,�!��9]]��K�B2;��ǎs-��U��K���^����^á�Z�ڐ��Ax�
(��e�i�a�o��M(����9�s�dt�o���c^��p��U���hO"�P5�������a&�.�̶W%��Jl�.O�m�9~��~)���"l��J4��~�,���w_����'FPc�0������](�d��93h�Jh.&��0�l�o�Z͠C�~��pdT��4����93NM�
"d���+�x�*�ϊ�D��T����@S������%M���5�1{uy�Ы��$'?ԧVy�⿄�)�ڕF��eK��6��G�S0�'&�qm�2���	����U��b
x��n�(L����	�	���>ӕ2��fFǭS�0v*�t1�u���Z�ϐlں�")��l~9'�ܻ�ؑ���AG�b�>��/jtt�;v�g�b�W�n��ܒ�B=t��g{�6lJ���ک�M+ǜ����xCV��|����DD�b��hM��'�/P�p��ґ��6�Ma��뤂)����Q��N�XH�[i٘q�?��y�?�~�)�l�bZg�_`�����X1V��B��H;[r#�<Đ�&���T�<00Z�o�6q��ݎU�����ٿ�HHR��g� �x5�2|g��%6l	4M���P�E*!8��2X��wͶ1���i�¾�'qGК����5�=4�Ӭ�M�mf,ΒMh���PEv���ge�$3�L�p���5d]qV."�
I�4�����T������>��� �$5��#�G���}ţe�ftD6����yم��;����5M\S�~2�Lxq�BZ�6����җ軟�Kj"�,�T�P7�1*Xg����SU�����%4[��{�,��n�o�����U�8��B2�����,�//)mO�>�샯5B�M�H�_��:�����h��+��YJO9Q������&��$d�>(R����bpZj��a�y�	Fb�D�>�*ʃh�4+��sS<:�oĴ��E*d���fc"h��|f���8��t��\�_����2��o��F����>o0ҷ>p#d�$�֦|E�I^p2&� 0�Y��C�]�HkqC�p� [-����ڨ<z�>�0B�d���+y�+�u�T��&Ҷ��\��жE�<�����zܜL~��� }F��__Q�����	.�����<�dfC����9�9�5��~�f�8��KB�{.q@R)�(���u����e}��+�`NoNU���4Y4�c�L�W�(�q�EB�j�b�+��\���f�f�Qp1���dY��<Gf2-� 
�Z����>D�Q�#æ��c��Y��V�W�Q�qX�޹.ݢ�i��w�gO���Z��Ss/kvA���
��e#�'�I-�WIw9Q兎t���Pm�,ק�c���*�7�ð��6��L)��>����O�F�� �	�@�@�,l�	p ;���jw�����c���
;�ŋk����έ�|��Y�*Z������2�sgՉC���rsm�B��£G�yu�Jv��}�ȫ�'$	NO@J��N򿝫+T���ؒe�"��G�z��������0H���$V+xo�	��w6X9��eml|?}�jK��4$e�"�p�(Wϩ��s��Zt�ֵ�z�����Ҷ�LԞSg+Лk�>a�	e`�T��-�w��oUP�+�.��B��4�M�B&)O�!f�{B�
�Q�a���3o���<X�����r��Ot8���q���g䇌UA��� _�s�{އ	a�ү��H��09G�'e���)�֭mA8_�\%���������5sex@�3j�tт��w��<�u�y{�Zr��̆6#q�t�I*�����\��Q��N��ٷʠ��=fKდp�oL��A������`3`�s'|�O
�\��,K�A�P3N�@�#�E(��M.�.ED�l����Qz�E��a����+��j�� �?�8o�,:�R������mq ���(��������_�惏Օu
��G��G~ �X�c�� N��j���0��:Zz�Q3�E��}W��/��Q�%����V�m��'�ׄ�Ott:�<�+��3z�F�2� F��qE��s�ϐ0cN$����W'��~�ƺ��m|Þk�
������o�g���Uul��ҁb9dn;� ���vd# �*p����x5<q_�2�6�vj��-�n��B>.����,�kϱ�M ����� >S�[Z���I�����d�@婢 �G�=��[���"?m�4?�ba�L0h\��f�o�ABDȝ�`������Kb�˽����n[���l<������DV�LB�Kq	�D��S�Y���G��������g�e���$��Rn�-���&&AV����}����'�X��\��SƬw�`܆)���_Ŭ8Q������M�-�3�ӕh$8Ϳ����I��r]�����	.���<��V���<�*m�#�P[�yA��V�f�|���Q"�>���\f)���Ƶ��W0VC�i��<�!���܉�����/��\���R��ѣ8�AA(^ji�OJ_�7�>q ��;�{�a�V�Ɋ@^!,�zڤ=���ҹ7�C�!w�ȷ�e:'"��h#���or�I��i�"�D�l��a�}OO�<<��`��B������J�X�@�ȼM��b������A
�C8S���1�(+R�'��j�.ュ���?=����^v�e��!�Y4�b����x|/�[7:D�l�����R�=
"ta��[ʈH �Kc���sn?�~&މ=	�O��x��!���y-�h�b��u�.�8�9S�O�.I��^W��x������<���Kd��މ
���Fq�M>����Dw�鿟����d�I��jȻ�CMX�&mI$Q�<�H���`E3>�@�ؤ)X`�g���  7]�=ga�c�$lL}�?��ٹ�����|�&���]
ӎ���O��x�a�W6lJ!R�K���A�����x?�0!t=�w�t���3gFVw��'t5	h����v\r����-�x=���kLa�:L�l�s[�`��=�3��a�
��Z��h?'��!>�S�)���h+�g��*�8hniIJ����h��Xb�9f����؞<� ��*�.S���;�I��&��St�i��w���g����)�/���c��H�ʓjV�	K��N3�F�����]g��˂zbNX�<�/�	�ޖ(��rb���䣼���%���K�LbB�{�0P�>��f�K����/�miBj|i�ã?�H�̽�Gq�K^�w��w�
s��ɜ�P��C��#n���� ��T*��W����� </	˞��Ȼ��|#vE3�|Jnp]%�����9	)��BtR�n�2��{�B�q/'�w)s`�p�;��w:[e����v�p�����x<�\��v��1v�=$9��_+>yl:�0��ԯ5t��L ��Ӵ'��9�Kc*��-�)��!���M�2�eG�aM�V&~H$��jv9�]�����lB����h �ϛ�����7xQ���a���� c�53�~G�LT�f���7)?�ŵ��^��M���ɮ�r���M�!#=�7�\Z	]�ԺԤ�x���,xd�۬�ʊ�eO��4N60
��Ҕ�^��g�����$�ښP~��
DS+�h���HGy,��ѷ�6!#�k���d�Rwܧ2����Ƭ��,s��yu�/�|�����dv�>6��1Q��=a��.���7�\�[mM�ə�i�~�Gۏ��;!���GU�f����4�����)'>�Lvw�tX���U��ɼ�^��jKOD�<n�����l4L��K
�ΐ���^��*	Åi_0Cb�Ak���4�ȅ�m�����lï ��SLZ" �U�����Ϙ:aBK��?�#僕�X=	^u\�C��F����O�Yv�H�܅��4"C�V�H�s��캎\XӡC�C���a�b-���P��rI�F�%{x��h:Z�oF� ��E�GŔ��V�� e����Q��6�}���^�F(W"�WaN�Vb]�[�{���0O��J��9+�kԘ���2�I��0uu�߬7��m�"�3��[0i���9_<5�������s�i4Zn�S�3Z�w��iB���A
H�#�P��c���]>��z�l����;Q��0S옲:Ck}(@d��f�3�8��=�m�P�W)�Hhjd]���4a/!|�7%49�|X�c�Z��ڰ������l)�u�gF��gm2�������C7��o��{}ɯ�dn��&��C _ϓ�^[\����Od� ��<Nroi���;�K�����4Ǝ_ߛ�ёz��Z�2E�|�\ѣ����x`0<�L7��"%���bY����Ɨ�~@@MaL�,6}Ȫ�C����}�O|R�Q��k)��pOé������5��,q�)D3�a�a^�q�A�c���^}��!�үP�@/�O	�9��ވbh���gr^hfY���Ǟ2�h�f�a��)��9�w�}H|=��u5��q1X	��^�q,O��T��(���>gqĊ�u�UO��C���J���EC�Ǽ�
�oO�O��f����bY\�ݢ#b��n�B������avOe��� ��[����c� N5���*�|����<Q�3 �U
������z��[�J+���
΄�@�Kvfǈ?4�@��8"�`�F�hF�kk��&0���m�f�2�m�bkIG*�M�$\<�n��|�M+>ӂ���7�X �ԋ���G��ܯ������(=&e��z�r���@�r$i����"�?��ϮFMq(��F4��j�+9�C[u�|g ���PH�+��33g{W?��璴2|:�*��(0��85�?��/^��8��Q�q��^,��>�0�8��ޤovQ�Ǎ<}���[�^�4�ّJ�Vj<�1O�j���$�~L#��Z�c`�[�������E��ymoQ"��.���u�����Fۖ1���a�3||}�N\v���~�f��FQ�잰��ǒ��T`�{O�O-�-�I�� x�N�����ח���\�����yۏ.��?���- HJ��V[���QH��h}˟DG4Ac�����*KD���U_eNg�	�yx��z��lcZ��xb������@�ٜ*����>�����o�7f�������b����P�Y�	I"�S�=��~�����r�~�\�*"Ƌ�CYߌW�@�k
�.L�O[��d{�x��U�y�-��^�P�F$t�l&���j�ъ-K<!��CK��Uak�6&���"<d]�ȴ���bA��U�g�x�q���ԍ��a��I	$N
��D9�f��]4�͝����k�'��)����^��RY�&[��.��@����!ac��*��(���?&-q(E��CC�F+�NsA���_��ͼi��^'��Y�5{�G�n��#e'�[kNe��Y�Ѩ��[:U����}�Gõoٿ�+�߷;O0ŗgT�s�u�5�9\��0)BYZ�'fU���0��u�L]�pmz..��*�w��4��uxa��L��iw�~9�Б%�kr����Pr]��se�>.�,'�qQ��Z8���R�����.�����]�q7<
!���7n0*�2���[�ȃ+����a�apz�a�@�ЀRY�,o�������2��Y:i�WȺ��3a5_�6gn��"��I���rv��0��6���O�E.�R �/G���Ա�-RM��8Px�ä��;�v�˺JF�a��y9��mHp�m]�Q��{2����'��^7�'X6Nv1��m��t�1B�N�2��L5u��\������"���ӃGa���2��Jxl����~���)��kIlT���R:C���l����'.,|�6y���l��*ث��@~rx�F]�E�%��\u o�#o'2�S��p���+�����S�>�/�����⎏aX'��M��(�0���M(�c|7����K���q8�ͩ�kN��ە�R����2�ӷ��ZU���K��)sA���8�ԯ�mD��7��"}aɅx6ҒM��+�e�+��~س����W�Y���tV�����������.�I>���*��M��No��w�Kf����O`f��°�@ ����z��dp�v�V��+�P�<0�^3��~�e���^��MW��3ӹ��c�Zg�p��|:`���͠��-w���M�Y������N�����_�&�˧�l��k�u"��oIڅ�@��.�"�<�Q�����i���:��rLF��tK�|�&��r������;�(�� �5��o"�&V���V�%S8�"%��ej�O{�S\*����,YqnQ��:���t	!	�U�����+O;��Ѫ������8�J���<��QfZ��_'��b�Z`Y�	��h�(��t���	����!ws$�*��M�K��r��{��VZ'���V��z��Df�d�����8�]������� t�����(%�YP�yʡ<f���s¤*�{���`4�!F:��׉�^Z�\��)��n$�Wdm�����g���1wk�o|�VOŉ@��e�/��Ĵ�""iN���ڄL@fF�:�܅�v����S;$���XIg$2dC�h�>�q/Hۅ�*��B�O�!<�C�-��c2��Qs����9$	˩o�%��^��JCq��H8a�j��'�|�7l|�?u���2�m8h�ST�5	����|?E_-n�H���m�� �p��"��7DB�p�������	�D
ܱ̈́�ٯ�?`�7�O�]ۅ�v\qp(�.L��oՠ�Ch�?\�5P,���&4����Ѧ\x��i�E�<X,��!�६�,��H��p~a�|D�iV�MOPg�aq�dy�G�O~���n {�^c�{ݧ^��z��]�m
�(1�]�D���i�	ԍD��XC�F�ʱ8�/g- �Ԯ�c��
u��K'��4�$�3g��c\<c����"�ڵh	�q"=�#vP�t�% =�Ii�o"[�}��q��N�r�Rؒ+�|>v���.�3"�M�¨݅���;���x
��Y	Mr7Ef�������9	iS|{���W-�<n��
����5��^罃�@��~���;ٱ���wk�����cK�i�	;��h���+}�\�f���Q��	s��Xa��,�Υ�M0�m/�u�,0�	�?p��?�<����9C;k;�ѻ��@�W��P�'��cy��v����B�n�!f��d����7��Nz0�������W�AӀ㣬d�W?gAY��%��\��SH�ʋ{�v��v�)�#�` �	w��l/rzWn?�})���h%�#�85�[�=+6�p-��w	��*��d�}U�8���|E�k��ʨF�Q�6�[��E��7�S!d�L
Ĭ��|�>t��ڇLU<��KM�����c5����� ��uf�9[͉�B��߬!�'���\U��(��~߬ͳIe����Gx�L�\��0v�!��߭^��)�����.ˀ-7��&���HsV�lW�S�O��W���S�%��I��OX�*Jw����Q;�Z�C�U��p�μ���?+��C����(����e>E����%/�r>B�߫�^��#���ءg���a������ɓi�]��X���[W���������H	F�66�۴"]�(`sP����ͭJ���(O������+/Y��r��W��R��<��u�U�t%�o>aYV)޻ΏN� r�0s��G�n�sY���ҵ����VC-��@3���L���q"&a�1
��U!c�W��kL\�� ����z:���g�ZƮG`z�砑o���?ժ�6%�A�r_=���� ��8�GJp�,_�݅J�FG��Y:ɀNu/��<ah��=�b�����\�+-�T�<�Lf{��}�	�FWg��O9(=3�&�?��"�����'���[�Tx@�����gkg܅*���ʍ�	�S�:��W&�p����\��s�e��5�+Ab������ymk��[��$yR%R��ϒ����q1�2?4a��c�K[�����sd�k��T�wPE�U��gBz/�F�se��v���Zt���b�<@���g)��Zp,��WĐ����1��R`��4@��4�p��`�n'�5]PM}�b+�xܠ&7ѯ |k�l5 ��8G��sk�l��5V!� �@?�s���"� ����}����iܠ��~����ؠ�H��l�6W���#�<K��4n6K�F��
�᝜���o��G��M)oM�{��,}�*���ə[:��an�3�f{-�� 6N�`	�^�^*3��u��鹓���
��	=���O*�ˡ�?�G�ǃ˨�k�*Sт�D"knض��<�Dwn�\��%h�'�3���~%��1��a����O=v�4+ M���KhGG� ��I&�݆2�}��s��]��(Ϣ{sf`hCh�&�~�B�U��\�NiWS5Og"�w�(-���IŚ��+n��Wܲ_n"9���W�a��)�ֲ6���p����=�O�cK<�9,�F������������\����������8�8@���;���+"��A��Hv�D��;��3��4e!m���O��P�Pu���Ӭ9�՟��_�n�^oT�ѧ2^�}-��[�nC����#�W��,B�� QFW�ǟ2:��
��o�Y���{7�۰�H>	���b�nٕ_��!�E�_���E#��c�rZ�Mt�l4b5����r�%&y'7,�;ufI�l�~�g�V(�N�N���H���{b� $*���)*O�c�V5�U '�D��p�2ET�tE��ͼ*8҆�N��#���̯b��qT�"�H+�C�FFhc�8�C"�<�$�l�qDo(����4]��3����/�(�"E���������c���kw\H��ci�:^{3*iQ�W]%dD�;-����l3��b��)��֪���k���/'J�ɯ�%��N�`n�[�3\P�h[�n�U�=X�Y��EV[ؖ<�!�|��Kܿ��݉M��Gh���cU�6e�r+�߹
�1Vrss�Զ�����7?#�k�I�����ۨ,27`�S��B8f(zF�{P_�<k�!}I���05ȗZ���Q�j��Fx�/K�	���B*�߱�:0����G5�}�������H�я~�jE���ܲm0ū_���l�Z�H��O�s�"R������vn�k�+ܢ�,��~̛����0N�4P Ǡ��sV�l��E��o���b��T �Bi&"�l�߭��!��eݚ��-�]�o�~�}m��T�_q�Yq�w@pv˅�B��ش�B�L�/xQ��¡��=-q"�j�vm�=��03Ty�b1�g����^�~C�gQKrh��'���}o�K:=F(�I�蠹�����`�2�X85��N�ܚR�H;Յ77Ț>>��v���]��;���d�vDW��'|$�k��B0����䷁ǭU��W
*n+�3-�M/ �AT:-	���h��/�i^KD��(3P�e`��%�nDl����T��v��hqN9k��Ɩ*61��l֪zC�'V��;��ݽ9'[�O�c�<00t��d&�1�z^z?��a���SfU��9}1m�IP���SQ�yt�Y剜s�$v��;�s�R���J��z��{J�fSڹXߜn�ʲ��#+�2�&���1�_��׌�v���� wӸ�K�C��	�S
��j��F��hc����8\��B�z�GAM�Y�tqj���~˕�i�a<��5Q�o�-�~b������/����w��݅� ��43�^�����zp�L����=��yԹZe��~pD��ܪ��ܻ���I�/��z���ߕ�s���n��뇺��u�J���#k��,�Q-G�OHl�f�X�%r�Z_�H�P�¿�7 FShx;���/5�� *�%5��ey��{�/���_?��R#��*!�C*� L�g�7T˕F��΄6�ь����G7��<��Rr�t����/\���\�_��4A��O�U��_?7���kګ'�GJ�q)K�#��h7}V����عc���:�a�T*�_ja��EJ���SG"U;Whz���?�@���q�!�(�X��G]+t���ֲ��#}F�eg"���r< �|�O�9�q��|e�;?�� +��q��hK��$��5����'4e�����_ũ�]�m��������R�����&4�����Zmq1�QDQ\	��@�n��F��,��\�D��S��<3����l�m��0�А�Sb�&��ʪC�Y��T�u���c��R`M; �.�����ԝbϗ�И�w���U�HO�Aի�3K��t�� ��q�'�L��kC�;�%T��݊bb���L���y�)巘�� #9����y�X���{��'�D-���ޤV�86���NF_�U����y�=	�
I`e�I�(zA�H��k�^��xk��7N�ũ��տ�ޒʕ����t&Ck��P�#����G5Dt�Y&9ƶ���ВN8���,7G	��x�fB�*T�;�-��,�# �`�x���X�o-���P�1�駇�����D�AΓ�d�a*%�4����������	��$Zoqπ�4Ӵ��q�.3L�u7F���*i�vE�������lP�H��gp���wG����#��	S�>���Nxw��'�=�����)����J~&��"�9���o�%�_qb��8�H�R�Vx�3��j�Omsh���/���?��y�?��"��$w�=��)�L5'�d�i�\��t	�I�����Źp��5�/ʖ�md6��cB�r
D��-rj��Ǣ^��_!��b���X�Q�<K�ĕ�
��^F�ٝH��� ���_W�Lk*���n-r����̝���bv�k>��$� �F��b���Q����&�лH�&��'���S�9ңTu��SXˀ��T��s���_h�ݺ }`������F6�Rqݕ����bH5�y�Mk����2,|Zo�����}L�33t=L0���ᶾ��ƨ��4�G�+SF:�I�wYWy�v�8���=;NF��2*f�B�G_I���*�����Z�:.xa�K傢ǜ�p�����X��<P+���
b_݃x.�ȑd[�7�h]iˈ����E8o��Mf�ɍ	���񀵘�xF�t��hb�#���9(ɝܧnu��B_��lGyԽFX���=�d¶���$#��]X�-�=Z��Ʌ�\�H�Z��:��^4b����s# �y)��u�+g���2V����y!��p�)31-b�)
�*M.��>c|A;�P��0�;�!���"��P$Cc2όʒ��-�׬f����d��J�z��73w���G�:����&O�Jiˡ˂M�3т�ߥy�;h������s[���Sڥ����	���h�ΔZ�5K���W�#�&��*i
�P`1�v.i �F��)��zPG:� ��� �ԙ�8 �W]�,�Ka���<��mR��G�{��kmR�`�&H�Pw����I���W:9Ǖ��L=tշ˪�{�z��{�np0�C;����ZL���&�'�|�Wi�dM�mf�;>�"+���C�⋉XUz��ԇ6�G�������'��a_�sU��GU�������	�rB(b����u����?�y�T�W;ȬUw�^_�,��;���7���WCnwÜ����U�f�q�}�z��T�Ŗ��RĦl�Q�V,�}��4�H���h��>TE~(�R��+��eX�TX���>�7��H8�h��l�<#'N<ܨ��eAO��K>ٽi@��}�g�gD �����ؾE�zޱ�����~�x�a0��nd 1n�K�� K.�� !#�%'ۧ��������-�lPv�w�	�$7��"�fsԲ��߀cfL]`>-�5l���T,�+ a�5��seRx��\?If'ʇz�i����?z-s�n�*�c��� ي-5���� i��ϵK�T*:�8i����Zk4B�{|ͤچ�ŴW#�r2��KtgL'��f�4�=���yL�r���Wѡ�IKH,}���A�U_��MLPm�c���	��\�F=4�f���t��A�u\p�Px�Q�E_+��!b�XO��M*	.@�����)~����U���8�gu!ZXI��k�z�)ð�r5I��k�i<�#c�8o�Q0=� WѠ��s�(�i���F�R�4���Q�o�����-��|N�ĉ�}�)�`��R��u_ u xf�T�F�k��Jc�Y�pB��e�:���Cp��r���596<ȯ�r�M^D��m�Q��{ITߙ*������kp��#9!3/-�5��Mj,)�wΚ��J��I�')a9�<� �e��ue@<�X�cny�"'�h���X����&�@Ms�e�]�/�I������Q�����@X��
�su�� AGzs�|?i��Q�b��F`r��8����Uo<��/R�w�f�z�oj�	̗l?g$d�Y!��}�E�@�of�����?�H,mk�eT:� �a/=v�Tޅ�麳�AS���ȡ�]�thB�T�o�Wj��tZ��44�c�+p�o;!$�ڳ��6�ꉓ�� �Q��D��-1򾖮�֥?[歐g�(ާx�,�������A�ZU��X�Џ�D
�_��Ǚy�#sx��W��)s�+�
��th�b	�&n}��T�{P���R�qX��D���N��	v�s·�ă��b�;���z�o���B]L���;�D�#?��z�����L��D�U�@4<0$�� �`���hlv.Q#.Eŗf���a;5���4�<8�	����8w�WA�c�e�c �/r���>�
��_��b0���6��몐��HpYO%�r�5Z�(��M��?���{���h��5�@�'a?D�/��ʝ0\eo���(�)o�]䁢���{u����������FJ�ߝ�G 0kDW<�z|�v�޹��W�n0>sx����%O��J�*Ei�W�KJ{����`ޛ�_2�YQ� �v��5M���PQ??H��ip�#��}w���Dղ��wuK���� �g�-�?d�s=i��^8��k\Њ]X���"� N��N�6����<�-�C
��cI��p+������uLͷ\��I��^Y��'t�$�zh���w~�c�	��UBA/��@�R.�󅆶`̀ľ�*���bc�{��\���G���;@/P#�6Gw��:Ϣ�.i��2���ȟ�R�!ᓎm�o��1�n`�v"7f�X2wO��o o�"�|�՜�U�����
�8��ͅ����nz�]'��@D@��c4!U�i��ᙚ��l�e!f���S���4(k��M�T!p%H��K���b�X����<�v��Fy��l���fS;&b|Op�9��Y �.~���^ivHܡ�D��y�A\�;[$�	u�	
ˋ����T��J�*0���{n��C)r���j�N6(����H���so��W�4��p!�\��K�A��q�>��D�[vt=�@�����"���G� kH�k��X/�j�:��q��
� �"�G������m�~����}7��W���"Fp|��ViRW�c'W������jҡ�3 
��G��@�U��O3����o�D��t.Ș�2N��5k�pOi!���Ŏ���&hE(9��LD�-F�������s���������h���P��V�lA��S-j]wZ�j`tA�ף!·���QjwH��� �C�B.��}nT���*q$]�o�φ�"����;G�%��o��o��s�5AY����W�� �U��ǎ<��d��=���?�fVnw?;��=*�/����?���p5�i����cMYSv�Av1$�z�m�p�-m[��b��m��v�(i�q[�%p���0)� �-�P��O�=W�K�+�8�$��Tp��q��ե=����$�:*o�$l��6�lٖY���VT-3�v�X)�5����pPM�>s5��dP+!_�ܯ*VL��::�&�1�v;��x�P�n��e�����M=�*��')7 4�e/�|Ni�"��6��9 �¯�7Oq����Y8��:�k�@E���k�9$M�߫��4
�_��)c����|�9�����`�l�*5��-ag��e� �����iR������K^�å��Ft������>�"�"��Qr�� a�Aه�r�SO���Crc�Şv���ʬ�a�<�+�܄f��t��D�#n���UKq�ʧ�&d�_C�Zf��U�&��S�r�V��;�}�kL1��Pt�}<o�gK@��*�k&R2W��3�PcA�s����b�1(�U�� �U�5���[<7�hv+�����_��+��|u:G�,��-85髝�Ekj��Ŋ"�Ս�Я�DL�P˙�z�R��@���P�����ym��4�_͙��r����]H�ٱ9*�Rf��z��6}���--���X�E�ϙ�X_��1�w��+l��$'=>X��&Z8�
�L��/x�W�@�U����c����v�����I�tӅ��pU�i��Ŀ�T����`=�KM6g�L�s�*iu�!9�%��I܏E����v�_]�y2] �,�h;�$�x��k����]��>lˬ>}�,�r@��ɸ��T����rr�����Ҥ��*�5�"��G�yž�7����y���̍ݢ��\��c��l���[���&�/�80��̈rk$����E"�Om���������D@,r�[\�ų��C�O�y��K� �~n�[]���ڥc���:����
*�Up9��Y&��'��1Nޭ��^[�������M	�]�C�~n�TI��oi��d�8*�˸?�g̊��J��R]=���������G�͒4����M-��u�jj}�*".����`�PH��fi�z��(�����o�D��m>dj�b�(�e~�J��_�k(�Nض��a�*�~?�o�XHhҰ�֭?��Z�hoaF[5�A>�j��	��H�^,l����YR�Q�ȿ�,�̘��S�C�]!f�^��xňZɒ�k6
8��]So��I�� ����S^)<DK�f�K��7����o�/&R��%~��/���B�2;=���{Ƞ�sk�ߖ��=݌�-<F����4������[�WO���JR�$e�K|���k)�}���_�	Z-��*��3�P�K�VL�]�"r�OZa�M��ܲ�{~��u�Kz�?���!�����A>�WW!�(��Z��/�,�u��t����Cz������2[rX@��]c����m8�}�?^}e$���mi1|t9���Ea�+��~1&��n�&9,���@��a��%�` ڕ�.���P�j����J��t�q��sfI�(�K[i�D����BNb�}��Β�^0�	m��֢%�yQ����#,�����̀/�R�=~����Ǽ��A��?k"�U��J����\Xrm`˪4������ߢ�g���D=�x"���('��CFulnK/�7$q�GWh̋X��4�B���J������A�m7��9��<�H
���6�%�f3�.vBe��f2ڒ�7�祉5^K��X\t�|���#�.��7o�ֵ���3�6Zo�ӄ���'�� B��e�PQ�z��	p�q�1�-@�hF-����=��v��4K�� ͱ'圜$e��w�tvJ�2z��g�V/��`�i���l�M��P��gRTf�]u<m��o���#ք[ˋ�>��=�,�$�Gwb��S+��紤�����1YW��y���wQVt74>Z�iJ3��X0��� 䡁2b�c��g-\����:��@L�̹U��)��h�y�EgB\�y���]�QyģoTcG��M���[������g�7�1�[H��,몒�m(��wb�� �4���tp��7�4`6�[&�i�Ҁ=�N�}�������@$W ;�:�Je�ُe�W e��-):�$.�";5<� [���lF`��XAbX�;�����+;1�Z��:��ku�H/b���k�Dh��,���+$��'����M�%�6:��g����tM�4VDê�m��A5g���f�D�>B�����Z�{jT)��e�1�'/�g}��o�c��5��<�X�B������u����x�Ң#,�����;�Q���xea�+}- 諳�g��.�q3�����V!�	��t�t�5B�ty(d*.6kQ�1 S֖e�l�z0�[��ז�lF�<,v�	�cl��͕���"6���;A�r9�+�.Y�gK�n�$���7�n��W�gk�N��������T�c�'U2�)�[:��$�	��گtc�_rlb1�����B�9�2#�a�w{�
��H�Ҏ����� 
h�X@dG��J�CR1�s�����G���eq�\+�Ys���J?�7��'�J�`"<�$�_|�]�_��l=��~�������G&�0���	Q��S��׶���҄'So֠��K�&M>�dRKoB��U�iݨ��\\/0b��P*�vD��a�tÓ��Fg�1��������݋�.���!v*�cK<%�(����R��$��}n��,�d�Ѐ�K��C��6�I����k���PD�Ѥ�c�7W�թ�Ǒ4K�B�+mS�����KaeǶ�`��js�R��<�տ�B�RS�:|�~-�9'�T�A�\�e�W���ƲK�ݿTkm.�)�$U{�m��b }/��E�q�V�{�܊��?^�]�Vd�%z��MJ>��^�'o�PA��Fo�S���&x�Ɨ%�G֑�yd���f^��sL-dظ�DzaU�xJg3�Xgd:��\�y� t>�K��_I�=0��a��<@į�*L�r��T?�Ȗ�a�������bs�:LS��n�tL�8j�ڒ�v"����b�vr@W�>'�2Y3O�c?sR�b��yMNպD���px��T��g�����i^pU�>J2MN��]F����l8�O�σ�P�Z�	�E !#Dt�?�pm]d�X*��Q��4z�)}��V�R��`=Ɲ�}�!ߩҙֆH��B8n��H;��PgCY�êl
S���0Lӌ,5x���@O�n��-�5E�i�x�i��gF�D��^��V@T��[FB�AJ���t�}=�FLX�O�����-8B��*p�=�<�^�w��r�ӯ5���Aŉ�n�?'�R?[��iw@�<(ҿ��B�F�:��QkZ�3�4iQ�m�%M�S��F���\0`�~�1���w z'G�|�g-.TL�3m'r���&�HnDKw���n�P\�����W�j�����h���H�y:�=��ڜ:�L�:X��\(��Q����YV�_�����%F������d���!��}R����->��1��w�<�i� ��8.���P~��m�TK�@�����T�(�5*kB<z,��
W����t\/_	 1�V���DmZ0��iON��#G�E�wM�����¢ht^�,4�|��v�ף��2�i��IGa��Ԗ�d h�M1�H�a��'~�A|K��=<���Z����?5I����fD�]�Xոj�3�:��ِ"� �qJ���O��U0���Z�Cķr$P�[b��i٭nT(�f`�w	�a����J}AU��qk6��j"������/���^�m$�o3�h����D�5��IoiM,�&�4���6S�E{kg3�o��?)�]���d��'�U����O���Y�j�Xq�O�/�EВV�~�3}�ŵ�����0d��m͞� ���5��˕˅�RN�tۭk#�'�ȯNۂٽ��Ns�B�����@u0�k�d��evMX����s��)��gQ��o�+�(�=���8a䴹"3�S^oG��G�y���`�!��x���J<I��[g�"�O�t���_5�=�5+��)��4�'�)� h�c�O�� ��H����ED�wr��O��8<T�#BCW�;?aL��
.	�`[�M4���P� ����-�I&J�Xx�����eˤ4�IJ/���1�t5n�ҩ�|��WHɷӘ��4~|�����T
�9m�X��zr&�? T���ʀ�?�������#S�KḒ������8{�ԩ��J;�O���M���=�V9,Є�ɘ\��57:�b��Ϝ�N45a��H|��ѯ�����L؟�(�@�=�T&(�z�v��_���Tm��4���*��plҦ����c/���{��8���x抗ȇ	��#�`�G<����U���R'a��� 'pB�e`���ߙ�I��)D5�����:����������"})�T�NV����]��F(�C�C_�G?P�;n���sN��T-���Sk�0��<��E��^=Ĥ(�kv��}��X��j���`�	
VG3�$%)���J'���08_�(}��<�$�P���<��W�o�O�j>Y��	��ܕ��uX�����z���w�h��~��4�8���8�c��'�����P�����\���0*��铯�W��Z�� �jHОA��6�w?�?�rB?I-� V����R����46��[�����M��
~���g��o8���&�m'<>wy��u��B�0�>��Ӯh9�*�Ʌ��i��~�MRN����SrD�G2�y�~/��a\�E�bTw�-fS_I�ھ��Ma	dZ�~8�f5N̔����"`.��;�,ž流L$����:{��h�^�׽��Zmb���2�#��x��Љ-w��SU%�+:4b/�*��yY�0�l��2QM��"�������N�6�
"���ShEv��++��@a3a@��^yF�v�α�H�-2(����d�Nq=4��2Չi T��c�-'-���|U#	���i�FI#�z��F7Q��'m蛣�g�'3w-�;Z,/Uci�\*H�c����Ļʖ�ߴF��?���Y�p�)B�-���wQ������pA%=Ҩ����=9���E�j�q��jњm�p���ֹ�������Gp�x��A��T��l�"�_�� �֧�R�1��0u���]�k�v��f����"��|}2���~��}�<�AR��ǒgΏ���G�\@5u�DD1��{�N	gMBA�B.Q��U"j	��B1�{�n��-8g�s7kc�Ut�b[j5e�@¦c�fJ�n��#�����}�|��hI��/��	4����Æ�A�tK�=Wgdʸ�D��p���&Q��m-?�n"q��N��Z'w[h��Z��9Fc�XQ��2?>��u�J�� �B�/@����;��qx.L"��Y^	@G�I�J��� L؎�1��"q�TnW�ܒ����k��#�i���N�%�d-�*�,��w��>o���'~rc��)PgE��VyS���Rz���0�"+��I�.�q�����z�գ`B��&H�n�ӄ���d�<\��nT�b՚d�"��\�/�� �A�g�ӄ��M��(�!�Nr�	�e�g�{�_���A:~i���x�f��QgE}Gg������p�s��SY�фާx�B��V��T4޴|g��=`S �i��'�&!s����Fi�p߳�n���g�~/��Ɉ���G�T��R��A\5ΐ��t�����j��������m[4��ՔD�+�'��S����>B�<�BU�4��l�j] M���e���bM�oӜ��&�LW0����g�K���DZ���K����x�Pk��xl���pF"��Fb�n �aI�����(�<	 [D���+ ���x��!�k�˃z"��R��0(x��el-���Fh��4��_��{��2�sӄb�Qg�8�)1�N��zqu��o���I���2Q
�tP���;y	D���'��f�"-�E��{,��L)�l�=|-��r�[�.��*L�}};1��1�Yk��䃏G�\��Y�9�%\�\~io@_/cs,}ⓣ�O�&�0/�$�d,���b.`mݦD�z#�-�ws{�����0�q�H$�:�T.���]���4���+e�|�5���9ILK0gw��:Q�}sjfH�nj�޾ǫ��E�aѠw��i��_�g��}��Q>�� �ó�GF� ��Å��m����T�����ن4���(ˈ��=����h������:��0J �2�˗{��Y:���!��ڴ�V8��jd����"�������Jߗ�S1'��?���ȝfZ���YP�ä501f�=u��7ca�2"����ܜ�8��Ϫ��غס� �'��P��T�o	�����Cgrn���۰��Z� -�gRl0.�E���Ģ���h��PIe^d�'�T�[Ȓ��3��ꀲ�ӥ��RbIS��H�{9�&�4DA��9�͂o۾�����G�/��e�I��&}�K|���0 �s�k�࣍3�`A+`B탕:� �Z1~>9RY�����5s��#'��|.&=Tj_��*�H;�ǡ�Zj��v�_X��k�ʩĜ����c2q`���;���0��<�� |���O����@�ם��!/��h�$xIiE�2W]�H�@��˷�(r���aD��������.Eh���J� 
���R|c�X�����m�\1ܥN{I��ļVH1~4QG1�O�>�O��lǬ{��p���
�������3<��V���`����Nx��e�|	�X�1�b�=���<��ZE����*����=�A}�Q�p�C]c&�ā��W�w()�pL��!^�Rx���=R��9oP�퉒�|�اxU=�7�ˌT;�y֦���Lc�W���yPфe��d�z�/�C��1LpD���A����"�5[����[{�a��!���'�ǟI�{2c3����\�Y�q�ɂ�G�Z�x,S0��C|1��wB����S��y�7�<&�(V!�:�%d�y4=�����$Ro
sqH����>R�NpK��`�&J1�5�s�O�����ф���R�U����V�ٺXx�KJ �TuS�4�X�U�I
q�BþI�����A�-����~2�����]�s���^���(�j��3?`�2�&� �S�l湻�$?��W>N3�=�\ދ-�ϴ��Ttf�+�>%+L�!���!��[� K�}6}��wq���Ԡ1u �}�i���W��v~h��/�x�Lk1�ϒ��\ڠ�O��C��C.'����
���	<\�@��t�Uqcp�9��l�����w���,4Y �Ɍas�la�d���&�����5mJv���#T��8���G�/h]�"�3"*x,�Ro_X!L����'�k���`�i\`{�ҋ�W��n�xPEۢ9+����k�8z�BY�� ��SeɈ�P�Cxv�%ͥ	�Ɍ��ĭ��	�#`���p���W�d�q��	��:)3d�*5z7�i��V9R���ׯ�8��c7�/�O��O�B���Z$Mz7��8����r־Ҷ��08*���������&l>�����撄�9U�C|��� Tb��Tն����%����5x�SV��V�۔��_��b*�v�ߝ� ���-M5� ��༎��P,X,��O5��&�ש�9�li�\K=�g��u�Ƞu|wH�v�!5�]����R���V�|��T�>��ie��r�	>p��qhj�3�N��BEΫ5P}\D}�$.�Jh�%7Hgp,���?;��+����w�pǪ3�/��ا�j�Uhk|%�1Z� 9�?<0>�;�11wn#�>�:�dY>����b�s߈�$}�V�E�M��c�K)�b�yD�onr-��y�7VP��BYJ��+����uyp����m9�D�܈e ��Ov��1X�/q���ݑJ֭+��P��FGҒc��n�0O:�HC�E��V���y�QS���RG?�Q���SG��x� Vt׻`]/�m��4)$���rc�W�Z�E�L\ue�h81
�*=����!'e�I���bw���A������嶋�3���u�+�1�X5���ufМ2L�dd:���&O��^$ǁ��:C��ȃ����Ƌ�4�<X��֫�U����\�;95w�Ԯ\ ���o�{��{A��M4w6L9ER?D�&P�߲2�"o �!L�&�2��t������G�r`#�'%nLҞ*V�9�7�Z��i�r�Z
�5�F�b��Z����#�!!��颒|�HM��x���}��7p��=��6Vnԁ�Ci)U/��3UD�{[;�ׇ��1Y��]���ɑG�L��%#i�Ӓ̧ҀH*���\����T&/���l(�����GAL��y���1�Iy��#����ۤB��U�!��x���.�f���8Ѽ�X,q����ě說`�1����;1O,Ή��2Ǳz�{��rb�R�Բ����7�Vi��	>W��mS�[x�Ϻ��f�˿��JQ�?8jޛ���m@F��x�@8Yw�1˗�(�ٌ<��g�s�i}g5�}�����9�5'h�fAI�Yg��QX�g/ ����XEuȤ���st�-J�ҠrONcd�Syf׷j��:P�����qMƠ������Xu:���������&tژ���� ��"�DG�t�Dun'��9�ª���T�~���K��|r�ҷ��O�o�1�n8�QY%"��&v~��yC�a�C�����[��+~�4��Uʺ5���[�Ӏ����}>��O��{�p�:s�>�I��fg���֥��G��?�}�	��d��o�n�d�y�J2%v�j�U��a� ����{ڌ8i�{�@O�;J���X@?��'i��Mv���FQ���8�m#7�	 HZ#d��/�v]2�����alq�;�f+b(�����"&�8�vbM+�-wJ��(9'�� �l��	-���0�<�my��8H��ϑ�&lm�p�<-�4����3L(��|��DxH��1�g�������(����Z*LS�8��7A2��=_4�г��^��M$��s|.����l��U�RQ��Y�E $��Z���'�e\:�}>�Q]���ő����>2!�Cp��cAt��j�B���{R��y��Xa� ]Bo�*�?%���������u���HP5{�x!�o	?1]�<��'ܵj sT����a�n�K{�qC�4u)+�[�n��{��N�'��K�l�\�tS�"��D�p����zn�\e�c��I��漡h���YѲ�@�vo@���`;kW!d-8�ק��o��H:�ǦL,w�rK�5�.�qW���Ĩ��>��xm^�Ժ#�o����wb����'F�$t�ܘ��`Nx�c��b�k80Qi�]����r�{��ZN4�[��L[�n1��9���(��
#�_�n��U@�y/3�ۊR�~a`%��i�B��ٴXj�"C~T�qZ�BCͥP���;�v��Zvm��}�����yx�؜l�#�-t(��֘kA��dא�`�8���<kJ2E�1�&%��B�� ��F)��^4�\T�[!>w�[:&����r}��5஽�O63���#9�%A�%��E�3����U6 �.���qàt����Z6�a0�@��P�^B��������A	)۸C�+���.�������|������q4b¿�:�s�A_Пq�˯�B�|K����yЫp�sPo�1��� ieF;�g�;D�kn���|;R�Ѝ�+&��QA��te���c�=
\�H�MjaU_3-��M#����w����H؀LW�8�Fc�y�f����wy�-��7h���o;����s0�]t-A_�6��O����o	q�6�*�*I��G�c�8�F/@S�5�)���(��3 O'g<���6�TBe�+�-e���E=��.�1_u_�V^��t�Kdo�X|���-��������/�j�8M�Ş��=���UEO)��{U�����nT���~�� �]�Q�b����ʏ����x!�Yͺ+�^�] �mA�Z����fmB��YW#}�,��^���B�����0�~u2�Κ�77�-0���X����ߠ�#�˙�l\MVK�H �/&T�:{��(��OL=v<���8S5�ӿ	h< ��\r�K�����3��	o�x����������O�+�0���+Ay<�M��B�.f��	�`z�H΅�
=x�[���榻��=���K�7���ھ6p��I� ���ǃD��afl�ajY!dg�I��?���Z�d�e�*���_$�BW�$�$�K��qH4��E�9�5)աl�{	�$R�Q�FX��q�����8�����g��J	���vXs����`����������k�9KP�,w��l*f7=Z�4������ZMV�ra�l�^Ԓ��x��!�<E��� p�b@�0k���t�屽$*
�!Q�pt����6f�~�*�q�{#�ȸ���8��Ve^|�X9�v.��m!O�� ŀ�x���* ���%�NERf��U/�J���-����0��k9�x|x�鿽���s��r4<�@'Rf�갈�Z�p�z{�pb�+}[���W)��<\њ�b'e�;Ļ����j�=�Ym;@����Cp�b�?�O�M,��[H��d�*.RZ{���v����yNbᣁ��� +����f�%X̎���U+����C�q@�Ǻ��a�q�����p���}l�1c���Py��*�|�G�*u����bB%x`t�w\X����P�G%|3�B$�˫�,�_bF��~�(ڹ�՞����Maw�Ghhz!�J5�tGs�y�^ZH$�=�
��'��z}:,�(���h(�V�'�J�';��p�Ne/@	N�H놭��~�b0SZ�v�}�/�t�n��#�~&)a~9�S e�l<f�:k8ZE��S{�f�į����	,�c,�l��W��z�?��I�Ʌ+��Li�X���@ǰ.A���gm/@�ހ�+p�n6Zڧ������w0\iWn~�H����RP���?�T
H[���9u����=-�t��a�9b� ���з��un�_�zfy���e)�i�%���w������5�;���!�>g\~dkC��n��{N7�9�GG<���靃6���D\!h��B#�m����>ۋ@@
ԡ�����U�ؚ��x ����~:�"��S�
[\k>̆��j�����2��pD`65w����Y������J�M}%9�3>s�p���j�>+�,L��M��	+��-u &Ay�iN��
�gld��ߨs�Ft�X��ٙ�ٞ�&; =�Ӏ�g�҆)�`O�xd����4�\��n7�N��~�NC�1!F���?���!���}�U��_7a˗�̯. �r�,<�Rc��Z
�F�Ғ��N����(]��0H��M��� J�@
��T�"�! JE_ �;�%�PpO�@ʚb&�K�Z�X�?�R7��/6J�)J��羴�Z�����(�ٳ>�"n����k.��`;��hK�~���v#�����8���M�s���_f�A�x1�%��]�����������|plK����je`o�*_��P�%�Ya�ձ��FR��ƾ�tb�&8�a@K���x\"���{ w�2�-����b}P7ϼK���t/�l�bmH"m��T����:p��eޑ,[�z�s��%3�YO�r��l��"�_��ʐl�kQX{za��ܬ�\.� R&.E�]��A��렂�Vp�.�ߐ?�=q�?�����i�vӚŇ�	�Ch�.��酌f��Q-�	�j���r�7��s�F����;W��1Lٌ�U6,�r���r?g��M%+*�G�PzB:g�D]]v�2.�.�b�o�w�uV�]ڠ��mdc�����)�_Ve������F���LKf�$����RO�K��)�=<Ӕ갮za�����ڭ�ozh'�w�S���l�����s�H����6���<?�{�Y>�r�V�ߝ "�n9���}T��_i�c�����9�G �̶�.����Q����8�[@�k��*�� C�<_ YȂ�m�=�
;_Y9�j	��3[�H��v��f�ߧ�����TP��4���l�n����M<y���TM�I#Bdl�2���|����S�N��N���,�6��̀��%�zG���0F?;�T�N���4�9��:|-T��R7r�>�'-w�Ew�N�w)���#8�/��!8 ٚ��UmO�n�Z6�6%�{�~�]�^�����!���2}E����*�)����Ҧ%l%]�m[-G��#����oF��q��"��e�8{��)��jyJ^������:+:ɗ�3V���
���wE#<��|%�G}d�+��|b���Y�C`��//+`��#;9�"yf��GpguP↦@�ĳ��H@B�Q\T.���2�w>�V۷�l�˷/�e�%�e1߀���4D�$� �[�uF�:w�-zV�h�G
��7	_m]^�w$�d:�ca��p¥���ZW[ ��-�&|��uD��)���rI{�6�;�!� ���Y�j�B� ��M{��s��OY���$"/\�駫�v��@�ư�V( �H�Wء8�n(�d�+ozBZ(n(��*�fvL��pg��ϔ�4s;6fh�� <��O��{�J5hW^w�F�c�Gw��yR�3�jڏF葃�ʶ��_h�z�س�����+B���
)2��C��k`�9�a'X婿��Z�;�%��G�r��Yk�������ן�4]�;oW���a���L{۳~��S�������a^ӄ���r�A� \X� ������e4I��)"��v�m$pϢ�C�����v��b�S5�j�k�j�mo������M]Ӹ�.+Ʃ�Q/���,��.��RʃTeP<UX���,��;@��(0�.?.jqUU�X��\�#�.��(������VR2�D�@�E��<���8���W������&��#��*kb	(�]������m�<�něbk��k}�'6��3�%w�Q�����en�c����UkU�����0axSh�i�v�9ff���mz�{%x����p�.�����~#��ӥ5��QQ�C�V4������d9I��4C�$�MQ���V+Wx<],��+Ӌ�eu�����,l>-�t��"�ҷ����T6\v�\}HmlX���ظ�S�`��uo�3�B$�t��Υ�0u�bC����{܂O?=J
���7���~�ݭ���m�;��T3F-i��W	�;��/�aQ�a<j��� �<T�9IK�3~CHi�k�(�/r�9���8����|���R�i�9�`�K˽0"!�n*4�['D��.T��?�l�"�j!kʞ���l�T�O2�2�.�at��,�W��!RW ����� jTj���~���/<|�M�ⓕ�x45I�D�� �&���˪z^�y�5�f�#[,�$_�r���c�N�C��jw����.%f�e�`_=��/ew\}�պR��Ǭ*����՟|׃�c8�6N��p��`�2lj�D&YH\����76mE�ɑ�\yh�{F��0u`�$�����������dj=i����R
k,Ns�j�F̢����<��1��`H~u8��zդ�XP����Jڙ�+-�hl��2h��Ѝ?�^���Y���Z��DDu���j�e��WkHD����C��IƈZ>Ee�9ɫ r
ka����3|�<���ʯ��i���u%K-���6=����3��NI���4�]ҫ�Cx\�q~��)l���؎m���i���b���j�w�Z�~˃�>�k�p�>�e�b��~7�F[�H���J��VO`� Sݭl��7�6o"���"�d��x��T�1�� l�y@���c�6�ȆZ�z�sb:��N-�פF
	èO�� 0���Su���j�A���5񀂕���ǩ�łe��k���c=�K�W�^��:�=�� r��0ӣY�m)k�#(7�!S�{`\�_wj��I)�i��ex�􎓲Gȭ�}�+7�I���L#�t�X�����awFd逧5y5ߞ�4b�?���c�f1W�S9㞣�,�X]ӗ�������zv�߳*��X�LE@��)��蓛��o��(x���|����Ʈ�6(u袩�?/��t�ƶ���6�fYt��?E}(ŕ�{6 sχT����J�|B� tRi�|)|;5�04njkT~��ʀ��v�A*��r_�ǎ#`Ǽs�]�Έ��.��Cp�24��$�J�˅�{X���q����r5�gaiP��3C��8?&(p��d�;v8=�3�>7��i���ADSl}bW�z�^�2�/Չ�0X���w/��H?���ł�d�������2D�` �^��&}Xݲ2�A�[t�j�h�<%Oh�M\�9E�R��c|�O���L�/�$��}���d�lM:�/ȴP�Dm�R��+�}��v(��ޜt����g ��Ҕ8g�����$i���B��K0
�3=R��V�N�O������iɄ=쳞MKA����!-��m ���z���g��!�8���Ė��%����f�*l��qr��$7��`0�����nG	~��Nɚ����r������\OMM뭗t-#.��?2(�p���>�Yu�����g!8χ�l��H�v%���p&����N5�C���!p	}4�����ƙ���ָ����e�f���oD>���iv��/{0=ѳ�����]��UX<m*����ˏ���)~^�W��JA`
���a$�L��Y�,4��*f�������U�y��Aӓ�8�3�|�+L�k����D�=i��%�о�K�E"��5H� C�@{G �)��
��T�]JP���z��M��x���QJX����bYr�T�R_)��1) �^{�JtS�V��E[�.�B�P�����μe�g91(.�k�_��@�{ES��3S�>������q1l�{�E@����\NɠF��Ho�����+�gke#	o���9nl�Ø(�Έ+P�F�A�q�Ý����r�$="�G40:���������$
/��OX+��|�yG� k8ᠦjj�P���9���=�?��A��;�A�y�@����Sи�=LJ��;���e���s�B-�fl3җu��,���D2�8�_�s��3Z��1�p4�T�(]-�>d<㊿�Z}@�\,�	�>�d=09qP��eJ�ﭕ�q��ʧ�}H@�l:����'��j�JY��6�����W�����-��� :|���a�����<���,m!<楓�`�o/$����9*��=����D ��mV,-͖�c����q�����w�7��'�[���PԄ���d(�m�Ւ����&�H<(�8���ܳ������u�*:�t�v&B�ZYݗeO��� ����dm-�����Tf/��V�>��ۈ�`�|*�'�D��3J���z4Z�j�4r�;*��lx���*�9�����iKpWY� ��'�6��Q�y9g���Wl��"�6�֯�TR�$m�L���'��p��P����D"(��c���ٍ�c�G�R�i�%�:\�ˑ{=��O4�@9O��~�m@W9��~����|��2Y�1n���;��?�p��;#��^��#:�~�N܊2��:|  ڀ�����oY�R%V��V�=E�F:�n�����v��c��#+d��l��4M�?���rz��Cm��9�D�Ǟ�T�<8�����Y��J�*yw�Zg�������@�e����={�޳��O��G��;�>��r�&,}���28ڎ2xqv;�%3[�l�)�1�'�T�.�Uo��=zc�h�-V���@�)Pe��i��".����ؤ��R\���������s�ҎLƩ�S��s��+\B�J\P�m݈� ��5V&��=�l��f&�0�Pݳ|m����g�੹� ��tϣ[莔m��[d@��@eɿ��\��B	�Eg����~!�� �<	���FD1 <O�Z`VϊJ�i�NOGX�;��@3����?�s�p�AQm��Y���8���'�HH�v�Ԃ~Ꭼ�hN@��-V�e���Oly0Vm\��������G���G����t8��u�����7��JB�*�O�����F�����`e����E8	?���S�Z�j��h�g��F�'p>�-�}��˒���R?ʂ���y��Dh5'p��C�,�Z9���V��p9����,�vP���φlGOu�F�u��?�����������%����Q����?\�����A��pf|q�_[�s������XӬ��ޥ��t�!Ѧ�p{�@�>Pv�O*U�+�=DFc4�>s�:���e3Yy�ƎI&5V{� n���Ʒ�VS;�Da����Gb`,�zXtH�o�����3I�O�0/vv�j;z���g��2�j�p��$~$�h���躐��r|"M�����v��Ò�ƶ�e;�땚cE9��
��y��� ����:qƁe����i����X�W,"ƅ�$ꑂ�Ѳ���<�@���k�S���i85D����z��|%�6��y�ubX-F�`�`Ǽ�<�n ��D�:��w�����dQ�B�_G��F�8�S9$��}�;�F{<�6�Ҷg�^�K,wg*lS��s<��w�
F�b���R�Y�l�4��}Ny�"S�ߖ����4�,$Z��.I��'��;������Щ��k��-�5��fY.4[a~���8��?��p�<�}�W���ioLi֮�+kᔕ������g�RW^�<��6u5�~R����Z�m��C�g����Q��#�W�	�GJ��Qpqk��[ә�ƧA�?ᶫ��]��o��HW�����,�� �Ƿ���p��=PD�a�&j'��"�Բ'E�۰ʡk(fʃ�?߫�|F(]���Q;�����F�xM8s�5{}�?�6J�"_��=j�{h�����w�&&[m	�I�`�R��ז� �3����Y+�u��	u�׶8_�
�t(�@�Ƅ�e���
k����A�Q��JS�P�#�?�O���Q�ng�� O���jɃn�^�a="x��,%�E��� ��F?�s�'7���8�\֡������2c�bج���|]gL���&Vk�@M���u%�JX}����	{��c�Y*ѮS@F�)��fm'{8k<%U2M��5M�����;c�~�|E��o���md.�@1I�&V!`	@ЎУ�۰�L�{آ�Z�kC��`Я.��.IL6s󱡯nuMo&�m�췫��Ua[?(oJv��f���2���2����a4� ht@�o�9��2~u�&n8,'@�)�
W{��3,mA�ɺ3����z/��w3�"]*m�|2e]:~Ʌ�
2<
�HЫ �ާ�������G��O���V>N�֌h�Qŉ��ʖv3Pł�ݠ�jFM2�Z���G*�kBn���0�/$�����S�j�ǵu��O��F����Pz�M�����S��ZJ����h�n�K	,�9������L����y{��
�T9���ߖ� "-�Y��fV�9�6����Q��rѳ��0�J�bޅ��Bu����5�󧈘�g��U�_wA����l$��K��DJrU��XqQ��t�`�a��Yn��d��͒��Yz����"L�>�u5wR���p/s���$+>��t�i7�^�3��h/���1XŁ6J��E��Ր�l���_t\�m�ҿl����Ӥp���J, #3լI'r�(�@��4�3-�=�*��]�{"�R��O�G�	�-�mo�٦I�U`�L��w���h�X�,��������,1���N�LO�hZ��8D�!��H�R�n.�P~�u�ljL��Џ���.�����UQꢗ�7��O �?��<�Ü{Q�hL�#h�J)��$�xg�վ�N<	;w�2�,��ՙ�����*�D�%�>�����5L��A�{$5�K^�������{H뒒�9BQ<�u�b��t�y��м����F1����l���E���� !����Ifٰ&p�φ��F���>'�g�b���໡�̣��A�5橦�/���W5L�V��}���'�1���l���wE!d�pR��,�iK�]�9����6�&�t��}@��N�c�M=p����u#�#.�r�%ʞ���h
�K��Y��?��a��b{"6�>c��2#BF�n���?�͵MdW��w��W��I�yW,�G`�_ c*��/�K���(�5p����OL�G��Y��XW[3 �]���:�54�j�di�6(Py��S��=���x̗)_���@���%>��p�P��w�a�<,�s��~��T�L�">("�<A����a��+x$�� �d�^�'UF&^�t������X�}�)7M�Ө�N��g]>cu!�'���j�z'V���p M�P��-r���v[��_HC����� <Y���i��;���c7iORe�U�* QƑ��	:L_��lK.�u�J�6h�<k�l�FU0"mAVս0Nl��p/��j�Q��pSO���Q���|�i���+w��#i)�&��-B�d��n��/g-0	j�;��5�:_�^X��ִl��Ntb� ')7��"�ށ�A�Ka]w���P�  \�*g	�O���\�P��Ts_�Զ�iF��:�-��-��S<CѺ�J��J���K��k,�t}�;�W4�?}�s9Z;'�g̕NL���4��h��?�1XN����ۥVS��
+��f9z�+N<h�q�I��4Á��u�4?�j����Z{����ി]- ̷suP��W��>ؘi~)T��wz�MY@�:�N�Lt�Á�ծ�h,M�E$A+)O�+ܦw�1��8�U�[V���hFp�C�e�3����/2�ŊV�gZ|�a$�#�D=Ṣ��0 mq��[�;�����PG79�q�������68�.T�y����Z�$p�q��G�������%)[*ɶۆ�~o&Hk����2�S^ ZW����I����X[Z�p4�}9Aec.�w�L0+5'pay�t��i�Q�;C��b���x���B��F�Lv�Z�J���HĖ�)Cä8��\Ai�#�χ��?!�lJA��v��XJ�����q��y;G%���#r���avN'yKB�l��>��nG�i���5��4;W �^�,m3�,񒋻��˭o�*(�}���S�1��)�#;,0����V��ܻ�N޹G�7w.E�Z�;dq���[��>9 ��\�۷����_���'bEv���dzH,�� �ߜA&��aU+�,�$�l����_���_�+�����4Qr\ʴT:�8�M
�L��T���t���86�(�IT�z�3s�,8��Fȵ�X	M����1����<�u������}-R]F�_]s)uTCh�a~l>��� v��މ �Z~�������uѓĦ�)~�sF*@��Ǝ(K��u�G���ʠ�`���_biAT�8}������r�-������Y��W�]��=�y��A3���А�kN��u06��RLb8�X�s5��'I:�5�D0����l_$X�D)Dt�-i�E�*�D��i���)-���I�}�ڣ�cH�����6cy�{vW������+�R�'���H�h;���3�`��<ҡ�E��faΆ�x[�_X1c�L�߻���`)]��m��54:��Nv��ǽ��!�}F�K�n� �{�w<'+b��/����m0ư�>��)d5���zt"��_��4q��{ȫ*���"�t���)�"]�%Y��|(�k���n�;�4�"��ݨ�95�E�.�i��>GA�淆_f�f�n萱^1�"��M%�d�{1)�{Ǡ�>��,�Br������4]�
I�����@4����f�a��]g��aQE�AfF�0t����~R��R��c#��]�:�YS{�6:�#w��q�G�;i[�[��	��^�fxFi�yI�Dsm	L�37H�.��]�H)��p�M���6`I�#�z�O*�����~�ە�d�'���m�r�a�ɘ�!���Q�+HgX�gs�����tk\����,�fH�[�$e/+`�0�x�H�<�D�����?��f�#��0n��UӚ%��.������\Nԕ�p��0-�(�Qte^.���l�q�b?u�����g��;?���ldK�z��*Zx��k�����o�u�i��H�č;���M ݹ�4]>>�`��V�S�&�����G�y��d(��(�a�0Rհ�v�V�'֗��Mx���"��]��p��L��r86�[�*Ļ��b{�I-ʤ�V~�qJ��mܽJ�q-�L�z}��1���]�f�|J�W
�0�>����Dą�K�`y�;\��n�������m#�xl��/���(�'@��M�E��������J� �d���?"��F����>Ej��Q �?'�F�ɸqG�#�] ��}�QW�����f|����Y ��I#�חb���&��/DVd#��z�-�D����T�Y$�ճ�����w
K�{_�p$$�?7:Zb�J7��l��:r�BA� s7��5��lS�T�������	� @�?3�\�ܮ;Io�MCݝ_�ïrb���P�xVYS���������8M�
(�"�)'>�Y����[�T������;��!�8'�IR>���v�(�b_�����ؿQ+_鴉�Q��5�>M�;H�s��x?c�ڀ�u9��;7��q�0�E����&����c�>suX�tGG$�JNL5�=�O7���A�c����� )�Գ��S�A�{�\��k̏W�j���~t�V=7�(#�u��Ƞ��z��������u�ķM����W̲ت�ƞ#�����)��Z��j�>'���s娗%�$�Nc�o<�O�
Ji���Z�:�������'�1��5�,w��W��/��o[DA&�Zpo����i�>���y az�:|.�f}�U'�c6�hP�9T��Q�C������8���d�.�w��<���,5�A�&�W�j(�p]���d�tY�R��߬���r�1�6��ŘӾo�͢_Rr'G�H�nnxʓ)��F��:| !m�46�{�$�*�aMw kf�Kǧ��B�B�^���2�Ls�@���?L�(�0�\^��+� ���Q].LgC���nO��K��H��beH�?Pb�%��}�'ֵ��	Ȓh��lu=%(�O@�Dy�L�E��,ubb�Z��)n�5�2c���b�y$������`5��]t��VXʓ�]}�\@,SD>%l`_�l��`[z˹N�P�9���w�u�����Ua����=
�ME�aeߡ�w#��D?y�g�	�a�D?�O����@��"|���U1ɐ��v������!�Rj8ʐ�Χ�ͨT>3�W�m�����l!�A��5�ڍ�`~����Qp�uJ����}��׵z`�!G�Z�@*��Xhu��y�T=��_kjO4p!���sf���_]!�����F^��Fمg�*��b_�Q=O�\�+Q sD�R��4�&����2��w��>w��{�˿�ȍ�x��jd&T.���2σ>\��.�<���5�W�Յș؃O/"Xk�a?���Q�7U*S��A�Z����̅���e`O񙈕�l�d�������8TZ���ER�d���;K]MS�G��2r�N�4Y4���K�Z�G�e����-_��9*U�;/����-�C�dȊ��q!�����ط=�����ȇik����ֽ@Y�3����$���K���5���w�	�)+�_'m�j	$�2y��7�X{������:ӥ��\�kK��!���H�sI\���9�ӌs�k��U���;-��ۅ=��]��u5(�8�@^�:؟ޝ架w�z��*��۝���S�h��K8�̭M��wq5�owr+`)��T�/ُ�w��)+�-��,?�<zbW�%;4环NcC}H0}�&���^�{G�96���Þ7717����N
<%x�<E����OV�x|��Sg��dfJR��7S%Rx:,z��x
��V;\�V�Ŭ�_O���\k(��o9��>a�4��b(�������!���uR4�2wd�'\\��u�l��?�R�muxO���A.V�8�H��qD8��9������p�#[�s�?>��!��T�ڝ����wVm'X�}M�a�iN�l�x,���kS�!\D��oO�g���R��ɱ.�e0P�X"L���nhH��Q��{<���*�m��5g
�|�~�W��t�4�qԲR��|_�8 M�1���I8U���E���1�KB}��(=g9y���zd�\��|5}�>C� k*Ĩئ�o�)���I�^��}�6F���@�^�߶؅�������aG	�oO��].g{��6�K��M�\��� �]__6A7^����[H�iZ�0�B]��L���C>���U� �\w}I��p�O��}06��A]K�2����н+x��-�7~�n��X'���pud%�`�h�3��3�Ԁ��s���_ �yp�Q�b�.��Y�H��7*�bGbX==lsW�UOo}�ҾƬ(:ܨ�?�@OyZ�8���I�Z�ԸoZ�M���ߜ�g�Ͼ#���fU<�,���݃�����?�����P�ɜ;���_��2a`q�A����͑���p��! �z �}b��qZ*<���#h��;�8b=�����T,���;���&�J�cv�e�ە��T�:�~��Rߟ�eΣ&�����y���㎉���[oo<2찰�є�s����y}�yVXy,�y8% Ҩ?F)D�+�� ���8R��,.�Rm�?s0H�M�U�o�G�d�C2oʞT��(b��2G*�s+U�_���a �r� qK�Q��8frH��7k$;e >N����a����+[�丐2'9�ƥ���u��o�RF�Y�j
�0�$���.F���%��' �3X-��?0_{9 P���,8c�>��@��qe�|h ��3
� ����6�]�dj��[��x7�l)Πz��*U��t�J2p0��c'X>7�X�T�j��8���E�+s+n��|?n�}����%%4�[Mḋ")C�ZJ�ۜŕ+����Z1�L� ��gu[��"�P�	����u��9u=N�k��0/�%�q����}W}"��wq͛��`����3���$#m�}?>;��ӗ���;�{^_����+����]�o�t���jtF���o�r&fL�n�z"��g���&[We���
a��Q'
�p~D.HU-+O�~c�^��X�z�5�K�]�:O)��I,t758�s�ٛ����u-���>)B�UՆ�Piѱv�����J�{&�-R���Z4���:����*�jz��s��.�q�ݓB� ������m� �C}����� r�r!|3j�`Cy&����D��L:�b�;q���k�Z�^�����M}w�9�}���Q��I7��a%߄̌��8�=�53��>4�E#�j�չb͇��@@��~n���K��)��9pD[B+	avZ1��З��#]|-�E}k
�j���,�Xx�a3�1
��~�� 钻F����>��cː�D~5C��.$22�2�B���>p��y�p��V�z�xGQ������٩��c�60t�p�Z�ʚQ`�,՗1#��4�.��P�ڀFoHqᇡ�9Ax��TLA��D4���e�E-A�#^d�5����DN�F�J�A��G[g���1�xe�iE�����lC9K�U0�/�H��v����o"���@5���@}�p���Z1��}v�ૺ���	�O0ӫ6�����R^g»x���ON�/�eh�ٯ�<
���#I��h^������~f��s�ɜ�̉Յ,A�#����&ӑo���<�]�f_'��"?�L�:%I��Ne����=[��K�X�ʽZ<��+�G��u�T����+���g�Y>�����)�;>{I�u�fܞ���;�q|�b�̜R�����(�l��ӫ�8a�E��S���:Jk�ֽ�z�~�T�Z���5] g��]?��a��C@<E��H�u7���7׭XP���(3���;�ߧ|3�B`r����#�E��(M���3IY(�ޙA=!O+��#O���3~F��pkΔ[,U����zƬa=*08@�z�U�0�h╁��v�(��4�Q
!b�}+f���K�?ߒ�� ��w�7}��w��O$��g���4K �W*�=�n�����t=I��!p��q�.��@ih��$i�L�|���,N{L��Ap�.�x�"d��_���9��kk��i��GI��l�fn�C�ͪy��=�EY�y��f�:�!={]L �.<��,�*L�Ĳ!�'D؉0�'���+��8H�R�x��;S�� ㇌�FKD�+�*��m9ykN�O�;S
�+01�n8�<�QA��Ҭף(0M�i�N�EV�]�zN�:����L�Z�>� �KC�=�&d�W7�`��t>Zc S���J���8Ňm5��U�ZP���s��C��E�\6��x�*]B�@^=�x��s�,��
3&n��v�c"��t����V�E��a�ス��y}��h�ޕ���t�7��kx��;'��#��o�k��_�a��@�>��IЊ"�T���J����<!����� �|�/�SÈ�ZN��[l���xO��^��8$2��k�8By>
-΃������V�9�$�a�y�=��G��k���И#.��=�b��ܑ1�8o�!�,\ �D������V���@|��@ME���VU��_��'*.�|��=�O�)��AeȁQd#�+��aX^�Q:3GGm�#�Mg�G�n������ RS6��{w�S#Ʈ�b&mºU4���"[�·�����jfO�4��y�(0�Ŷ�Jw'Ńl�pqV�M�څ�+��<�����l���M�!�X^�n�%YQ�_S��G��Y1��S���^J�U�����?l�n�9�:�hZ��'�~���&r%����Q���}S~ܟ\Pim��Ӭ
ñ�h-L4K��r�l�⿆u���U�b��nN^����>K+q��#p��]����P6�$����������.8>HnL����V�n�#�먻\�pK��iRX��e�^`��<>v�����h��b�{0����o����+��O>���_@�D�������|����!0�23�F2�g��r�!�g�ڞ�����q��`�d;��8m<������]"$�A�H��gD�ҡ9p��&5�G����U��9Ć�Æ�����[������JR��nH[�%��&�2����	�0W�-�����B�©!�[�F �W�����QM|��J��܎eI .V�
q@u��V�2�*��?�;��A�8��˾�Tf��a6u��E�a��)0i����B���l�J�1��ځ��2��ɶ��tG�Lଡ଼67�V����w�Y�ܗj�|��T=f�̉A@�Y&����j����(�#� (0ܫxF��]�r(�0/��3`B�ߓy����%ץf��ɚ�=P�wI<�ʂ�����Z�\@�{����ϕa����|��,����9�����7�|&a��]����e��E�ϛ-�x�k���W�G��$�#"�'��[����{S\t�E��=���9��Q�L�����U��JB4Q3]/�39Ed^k7��`\���HZ��Ox�{��i�C��M�^���O���|�RU�"[5$����%�"�P�a2�4����kҍ̂��+(A&(�#�(�Q�����b��c޳4��'/����#ԟ�2o��9R�&kâ[1���)�Ze H�6]k>��3��¿�L��-�9�%��MS�����H�z;��A��j��\���{�wZ��}�J~�U���ǦT�pI�{�i�ҡ/�Kb�V�@E3K`C�O)�
�,�^J�ʠOMǱ�}|��(�8�ƬՎ�S���޼^�������ev͒��Z�<C��h�0�C\,�ԣx��w_�o#[��`rC��X�d4U~�:�5�W�t�W�8�w��D6��~
�"�%>-A�4�?�eP2�*2� q��4�A'���T��G��;��{/�����Ǆ���u=� �:%�S~��.�2�2�X=���x�. �]ŊnM2��ërB��Q?����HH���~=ŵC($W�i��/�v՝t�fSS{M�-Ǭ��ޚ	��Jِ�����>��r�-P�<���<g��n'P���>��F<���m�3�pw~l5��lUu��c�{wPco�����-ٕ*��9h��ˬ�=���G:���[P��&(;燈;VYJ�Z:,�S.��?�Ϥ{s]�� ��@���-6%���sZ�:���a̝R�,a��������K
>��ױ4B��/i�$�F�'�s'zA���w�d��iꯎ�v�n��w|փTbD�����D����ؕH(�(��@��L:�na� � �i��`c�hɜnoCF8f;�URW�,k-*ąg�&�zo���y��tҮ�'I��;'a/�x�8���x8��n=��%,4�'�<�l]��щ�Ԩ�RN��x���ob�:�3���30��Dß|�#$<�=$�����:�И:��J�3��{�3����?�4^�/h1p�k�}��1m�YP���F��� �g�M=�T��&Q���x~*2��êjk�+��ҝ��-Tv��n5I�l{�V��#��\��L����W�2X@��<v4ȯ����dߵ�ݘ�Is>wLDŅ�OY�~�)lHϓ!Afq�1��\g�e�e��Y�?�����N:WU~�≮5��޹ZjşE>ЬE�!�WB2�`̪�	��i���a�K�������f q�)ါ��I9A����������־����PmO��U�f}� o���5K��� w2S��������o�н������"pB��g��.t	rjmI @ٽT,v����RA��Ԧ#w#~��i��ImA(y�C��;��¥�"%d�S�=}���N��MDv4�8$��o�1��m��?��'����0�1+f"ܺv�i����m�;��R�A����eh�>OT9�wa�?�%���(��]��QAT�tWwbL��b"Xy~+�Ն[˪��z�)���i���;�)����f��j�r���;Qr<��e)N�\o�D���O"71 ���l��Н<}��Pjy-��!��'Ül�n��/�r;��2��)Dl�	��o�oћ�K�{�7�=m�C��a��^?+�-ȯ��^�t�4�W_�{C'0�16���Y��Y�z�H��е���^�,^} Ad�]�D�v���#pH�6����d������\���������nW���C����l5�1�{Y�v9��^l�6�~ٺ���ňwNE(=�l�ߖYRѷnO�|ў�Jj���gӣ�N�;��ގwF��#s�]������/��m���ro��\�<���dGX1}ץ�o����\�������BZ���fވx��G$yn;��*9h�rtw��sC����
��x|�Jžų�I��C~�����3;���Ў�������ԫ�rR0(T�=	��o�t /�?$�-^�>��w>c��������V{�A���Ԣ#����%�<+O�!�� z��]���QPK��}�.�=�K�~�ʹ_Q�Bo�Ǯt����۬z�V��W�χ���:.M7S۔�����ߏ��1΄9خ�Rw|c�k�Ƞs<�@����}osT�-����܀���=���"$��+�axfYP��W�#�w�o�|bA�`8J������M��vU�v�w���NP�^h��XP�}Z��K��kT�?m�� 5FCR���X�(��I�󯁟�-�7p��4{��4g�$�c}k�i����٢�^��@:���J8uu3���8�i�o��8�G4��0�I����u��M���׾��FJj�r���bN��P�?�9ߍԫ��Kl���u'Q'�Nղ~w;�?��.��q��pd�%Q�bx�N����V������U�W<D��E���6���r;��ى/��ʟW�k��_te�z�@���D�����F�'2�۔~7�m?��Nm����@yy��LVb}��65��zl6n-�2>z)B��%7�ؕ}}�,��o�41� �9C���W�X �_U�<a�'3�G�\�X}R��o���I��'�>R��O�t�*�I.8tS�8�C���dg j�0,��mD}K�lK�5�V&f�{�u����k#֢��4�]6��#�'v�XEUg8x:��e�I�P��Y���j�F�q�ms�Dy~�쌦=+�r�z�+g����4�D�q�<Tg?�D��]]0"��J���K�,�>�}��)�|2Zm�S9����zŗ���l��+�:'r��^�;*�H
4�z[?KʙI	��dR��?7��@�*���稏�t�ѫ�5�D��~o�㷱F���4x̷u	�?���T
{���j
����H�ͤ�&�QA,̂�nh��"= P�Z�}��sNб���}���i؂��d�ܽi��X|
�,ņ}{��FUg�"A��bke����1�TA��R!=�������u�(	��=��i�� �^K,��N=Q��
K7j��������tl&%��증$�a�t&���a{^�[��e�KT^��@�����M"�_o�_{�/��ط������#=���o�c	0*��R�.��\i���G)��C��1���B���R���Z1py��K]�go?9_�B! ��?�������<�X
�R].�M�Lz�.�z�l8��v�砘$�Us��������ʏp�Q 9��R�������箼�P�ylM2	��_0q��N��	��C
�ԫ��p!��^)S����@��S:�Nu�'05�˔EB�$��1��U҇,1J���,ːw�������/�����ضh�-��$wkj�B���U@]*L�$B���1�a�ƥW����#h�95�#��/�,�u�+�>C����'C��dkү�tW��w���u�š�3g�ܣ��!���l�7����?ny���|�V�Q]��NF ��l.}9)���G�,�+�3b�����Di�ܸ���|�M3y]���02�J����YZ.t�t
��wPl�O�%�o�?�����D@w���HQ��YjJ��x��=PD�HH�u�a5ȫ�Eʦ�f��К)=[�A���k��'��?C������~pA�p��q �X�T������9�c���֑~H��т��"ٌ
�Y]ݡ�g���e���\���){]5��Om��#�~�a�:�yU�$��۪��^˱AG��~��Qi���������Q�,��n*L�W%��1	�4%�=�?� 7�$Yʵ���<6��
�
�ה�F�ŗۄ��-�Y-�^����HTrY���Uuv{h
T��G�>S�Pr�(b�㷙2�za��J���8��?D��ʞ���X�3p�w��)���zG��̙50s��"��&��w�c��x�M�<��uv���Ɨ��)W^B�o�F|�2�0�/��jbh���ٯ�P:&A�y�X{K�[��6��0	B��;1�V�3�7�05v8�1ƿ_�ѪPu�8D����wB��'�+jq�����~�ʐ	g|�X��ʿ����4%��t�\��o�"�f:d|�����@�dc�OUI�2��xS���XWf�!B���KJڟ���pQ�4�!\���5=7����m9n�!���N(,�����&�E#S���$&�`�(~\)б��j##��=^&�dfO�/K�"��\�̧rts�r*���c;|����]�ugm��%��dN`>H�o��<����+�Vy�7# &8��4.c" ��״�w�t�
���C�Tf�}��h�ٰ�<]Yj9u)�Sm�27Y�� �kq
r�摉�72 r���!�J�yh/��r�I���-�����c
3�[xW �N�N�)ľt��9�ކv2�g���U�(�W�:��2���:$��M�ڋG�hNxf��ix.�^5��m��L@�;�׏i�GIX�"����h�/(��J�v�zdAK��r4�X��,2P���S�/�zrE�H��k�ߋe���o��l�-��,pN!��]�a�\jiI����o.�@�x�.�w��z���Fy�!7�,G�H���焔Ш��3��d�T%�ݱ��d�D�^�m��H~b��ǊDeP�B�� (U\>��e�Q���W½u��+k��9���_֥dI��5(�/:�A7@a���A�vFnG̞�>!�<�����_*F��-�q�����b�WGs[���m��;:�}��s���P[��D~Լw�j��Ru>r<���@C2���W+�G2D|'�W ڲxN�ҧ�̶�=�~��m&s��	���������w�p�Z���c�AҖ�9�W��6�P�
���VM�ؘ�p`�T�Ew(�又k���2C�Q�G�����X�E�b�u�(���; �	��z�� ��э=W���/`�_U�DE�a{y���%.������ޏ�B-�,�Y��5gO��dG�)�����`��la,/����ˎ�'v-s�
����l>��J����X�yD��U@���d.�B�fι�P%�
���ȴ������)�h�\X�r0���p��9��=h����G���E�}#��!�·j��o��1�4N�4��ɣ�b�@��w�=&��"b M�a�@�#K��� �U[���Y��w56N����,��<w�apCC�3��}0�'�q�uZ���y��=)�@�离^���w��hi����`��S)������l�YXƊH{��j�ulC�t��/b/�Tud���8=��>3������I�9v|/%��]qE������*l����K�W��ʓ�/
e=�p��㤝�%D���hX1���{OJ�}�-8�lFuB�&m0w0��/��UW��j��ReO��͞��"���&�N��㚟_sIdN��#�}���uE0)�eb�U?�p��*�r��Y(��%�����c4�:(��R�g`��.��)X�����y�u�}F��<�?Z_ڤ���p�"���J*�؋<c��u<#;	�d�+�緣E
Q��x�"v���t!7@
�AW�̒���"%n�An� ���섗ݕ���zY�D~*�5���R�*��]�S8�"��P����)u� F[�ը���7�����YPJ��W�Оכ�E�QQ�.2�Rñ����S<͓����?+���l��=���-|�� �t0��AwɌ��Zj5�8�W��'����U�8���m�����2Z��4u��l�Ͻ�R��fN��+��g3Q�U�ɨ�으��.�x�Z�4��p�~~��:�"d���v�q5���m�x�'jR���(� rjH�o�Q3gk���<���2��	�"�e/N���emK������ڮ~��{������1-����:Qy��VN��>�YJ�F����5�XM��Ģ���IQ&u���-��9���&t�}�kWI��|����B �=�]������gw�g;�P��
8w��f,^W���;]ga�$�ty
)�{��7 �<���� �öly��!YM�U�5��L��q*麡	V[�'
�#v�Rw�d.τ�B��bs����ILZ+K����oN�8�Kf�� ��ߤ�_�6���#�����2�fww�`-�N9��8,
U�@�Sꀫ��4��W��Az����_�Ef\L,HR�KY�_k��+��4�_n����u�np/HO���2�p���6���K�'w^���Pˍ�coa���H��"�¬�a�C��{��|��r��e��M.�%PN��-0����g���q�ɳ`��K(�˱8DE�FmO�&vɈ�`5͸8�_\�W�3��Y;�(+�S �-�K��yrf��Qp�;v�z#?���D`=~�oL�+��`�5ǩc��R�L�;H2���0V4�T@��I�q!�H )wB�)����:�Q�b8�3��;lS$]�O�LXI�E\����B=�&�ȕ+*nqL9b��R7b\�{�qt�m �%���)�����Ea���V4}�K/�i�4�V��k�!PEasl��gd+:�$7� ������_<�;�W�ˎ��Rӡ�������"ז��[1�Idy�����`'�F�D� (ˤ��Hm��U���ܙʫ{�|Q�/>���dkִ[�qC�3#�<QxLR(>�)
7��9n��Ä���������e�Q���@���:�3���jv�j�н��Zh���cf��.-� �m��v����\^����Ƕ���0�)�fOr:E}�x�A�S�������Q\�\��J:?�Uم�U�yx���ݠo�츖�k�w�ܬ��񭔮���i��#ε]"FF'%��gYM)G����r�V�QL�E���"zM�H2Jڣg�����[GY�0kKf���7�-{��=�������a��O�R��s�D��Z�X�{d6ZW�g���
�_���QA*���9='�2G���Ib+�BN�I>S�f��9��l��`e����}��}8��_�D)~�f��$�l����%�(Q�n�:��7\S����Eyu��&}e�~���A�!�e�]�YL�N�1�����v�>��P�$�yf:iqW�$�w�>�\@�mC-q^j���}�/��E���t�py��߿�}[����ġD�j�P�6�۞�r�ӬEx�p�+�����'�����Fd�|�uBJd�4���	 �E`�ǇBK7T.��[C}|�+O���`j%��x���
K�a����J��*j���­ַBTB�{�Fr%�j4{�J� �)K�2)���x� ���yv��\�h�x�ej��	��9#�����RʘX�N�e������F��tB4�;��R �����O�Н��;�:D��5����tgNp��,?y���li����آ�|3�T(� �D�@�s~Y}�����NJ8OXw T{���}o1.i�.t��^�1�p��o�'��ށ��*�?��3�X?�Z�� 3�2&0�]��z�F.�5�����H�ya��g1
�|kk�'��T�B�9�Lb��H���,,�hnC90��p���vY����-�
oTݲ���w��l}I�ሬ�Ś����~�N��v���-ɘ�Qؙԗ켊�j	��â=�a����X�I)��,4��i��D,lb��TG�8�酻���S7(￮����D�iÁ����D>��E%4�qYc̚�����JK1,RZ�ɱS ���7�O��W������V�v��Z �|�^L ����0t��f�7��L�ك7z0�q>їbl1F�n�g�����R�¾�u]s����ݣ�U��Dң<�\���pߥۊ����MS̊e�	+����,��lXC\�,ȱa!�1�����������r�0Z���y��z��V$<�5�kyR���R ���6��~&3�@��=�wU6��p�/F?ǥ��ܝ��&>Jw�����7�o�-:)j�̆8��L�����2i��	�0���>�N���u!4��@+�^/����2c�h�gՐ4�c�ػM&*�|��?��ܻb22�K�0�h�Yp'�9��C�.�Q�0�D�9A?5��Fv�<�F�=E���rR��Ǣ�)��YP�%��NP�:Wf�n�y���Iq�L�\�\��6����Ѭ�T,�&A"��l������$�ˬY��W�T�$B`����r�$���5�+s���:��'��K��,�2���!�Nʝ���O�����ʯ�����eO�!� \�o����6��5����xͺ��\K����y�Qf�*�z%�;�9��/���ђD�;�����j|��!'t�|:޶�9".Ҍ�C�r�,gbl��RGhL�B$L.��k�L�����������r�tS���]�9��KX��j�T*}{fބ�{Ij���V>��qF��͛���j��^uP,�u"���u2��e�3�7�qv�l�iņR��[���@M�{/|Q\�����ԩK�)������Y�̽��d�.�<����"��Jr'b�ּ8�K��� �p���s��T�١�,�%jP�O�v[�#Bv� �&#�NGK:�%c�!�H�;</��ӬL�N[hAhQ손c�J�,��f���ޚ�~1:�� bʸ�,_�y�� &�XK�JUuA�B���]�1��S-s���K���҅7xqS96��%쩆Gg��·���>�Yŭ&l�b|�f����2ZHn���u��X���u�cX��&<1��|��"����H�h�+\�E�
k�xb;�B����ME^�P�0f$���2e����[����:�%?T���63�Ź��_2'�p�1x�/��N�(D��"��ו9��I�G�4�\�u�f������˓'�yhV�q�tF�!� ��_���z�h6�J=�{>�g8�Ele^�ߒ���u�ɈsP(��C_���ƽ��葿��<پ���#��w�x�C���CJ*h�V�^���.�Yr�1+�x㍣�0�f�i���je/A���9��<P.Q-E<:�W��o5��yăS��C	VQ:/h�l؜�G@x�CT����.��
G;!�ז�-_���=����l�L{h@�	�<��cSx^�'��{'T��"a�� ���tK�`���t�X 0��^Ɣ�G]#;�ݟ����S���h�g`�~�<y��m����ۚzX�p���Uhp�qf�2U���н������n�e�1�J�h�w�����(\����N%�`���%_���+R>��R���C?S��
E�^�܃1��M,�[U!�u�O��R�b�5R4�*��ǻ��!�ԙ����T���4VR>�g���ْ��GK�d�����ъ[_���Y�e��:�ρb]RY�	�']�~%[����C��4�Z�F��tw��ڪ�=�
�*��d/5e�5!5���Q���M����^�":�Zhd��DWP)�)�`<�IDs�A��cXӾ��{ݽ�H[&|"�eV3^ �*�SÑ��}�98����	mse����Cp��c+��Z�/����}˖��O�U�p5���8��� W�V/7��c)6č�&�m'n
	P57y�M_���~�q3Y�Q���g�ItiF����1� ���Yip�0������Eg#Z���wa}��w����t�X�D��H�� ��IE{��Z�^�rcި�9^&��@�?��6Z��Y/�8��  qA����9Oȏ�g���kW�].�~�%�4���|Gd�o�1�E��t/����b�w��Ă�z.��C���hꍙ�!	�.֩�`����aSO�qm9MY���j�9�T7g�R����BwQ�-l]~o�$w��=��ʂ�H������䡢�g~����E~�X%�x%Poz�:��-�O����ߓ�q��o����Ο͑v.;9 =mrOP	�f�g�(5�GU�\��ⲻ������4�1b���1m�u��B\����AL/���(�9]�D�M�t�صC�2x� R�8�w�E�Q��8�l*-5�����_��@��ݯ>�4�g>̀���C��zd��Dcҡ�T���T���an��ǋT{�ֺ��t�%zO�u��5;�j�+��6��� Ղ�����.2��A��;ZP�%oO��vppL\U�d�,� �~5H&	���&[��� �y�?���67�z}V�<Y�9Ф�֓�٠��]������Qx���G๛X΋X;���D����|0��#L�C�5� 2�@�X�LsN��gS��~d�Jq9����J�ɱ��ԧq�����V�8�J=lL�X�(��)��~��hu�u�$6�g-�H5Y��͇Fu �7]�HK���v�I���yR�p�\��,�������.M��ź��I`�:�}*��;�F�"j\�}�OD}�|t��CD��Q��,É�\=�Cq�rzm]�Ǉ�S�n��������&<YM�	Qc�f2	�h�3�=R1�gCά��]]Wr�9���n�׽���p	�B#�����ޟ��;�af��:X=_&g B��X�a��	����W�Yڂ�㠫Fʹ��T�g��*��T�a�9������IۆY�����d"�[g���z?x�fkK�p��p2>�Շ\b�w��,�6i!�j#�'oe�)���8o����ώg->��W��)~$��bJN�t-�bb�ߟX1_Y���ł��_�����io8 ��Jx��wo:eq"���#���8�ϔq���������C��c0�eJ���j��P�T�2Y�����w(�8��6�bQ��$����ʮ�д�{�[j�g�����ڪ�µ���q����E�lU��*���J�L$�iР�Qu<U��65���/ �WЄ��쯼
�ejd��T^gs%��K��h�3���0,��,4�v�S�X���d��:�X�は�$�'ጻ	��.���0���[�z`~�4�4ѩe�jz���.ѧ��K׊�~����D�!qL �)�YT'}��F=u��bU�4^1f�%{3���bk��=�·���*֍Ż���|��z$�� ���V���Y��>���Fnic�r�F'��+V���nm1&���Vn�Y��\f����q`�攫���]}�=���+���S��:6T�+L�k0޲��+8*�r헭�8���(0+�܆��|6r�� L�?7-<����� ��(fIլ�S�t����Q�W7ܪ�[8���|~�DfR���ދ�dh�,>��ւ�	'a��,6K8$XΜq�Z��;�Τ�ݢJqeTFkW��D:��g ���j��k���K����c}դ�0"���j��U�7[ܻĤ;�:z���,���`����&_��g-�jC��U�x�O���p}���.�9�݇���'�[���ރOu?�7n�;\�
��=2�5T�eoQ��Z[����1�W��u!�_��@�쵳��"*PmD;�.��k��%��c�0,<4�A������B����Φ3:�����>���}�\ē���{wש,,� ��Ֆ� rϿ룳`39I�~X8��*
1�Sx?٨����x.Q~O붬�zbH�`���e�ǻ������S��8��DӚ
?x/م��\3�DS�NÃ�l�c�����xv[����&�:@*F8��S�cU*�:X��h0N�#�-�.�F0|1�P;�J������-e4S�K��߷����.��%�V}[�f	����:O٪�����ZiUF��cԪ���h���r/�
,���5F���b}����cA2~yy�&U�fq��P�� ��14��i
UHjbF�,�u�b���+>Jx�
�ǂ��Q����%�L�7:YD�;��%�f��5n�*r%�O�	o��f���pF^7�[��'ծV�!^�Ua�.�{�I�Vgu�eD����
]�F�a��K!���a�d;6��yM(':<�#��9��h,\ i�He{RW�\�?�>R?�+�v�D�ᬚO['ۢ`|�4����کխ�`e/�]'j�2���hy����8�Td�;";չ�e�y���,t�y��S���پ*~
OpH$D_��-ZD���3}E��,<����2T���(�.�I���P%��h�#�A���^#Z#�\���i�J�:�X�:��~^�ADTj���9@�'NΜ33C�qN��O�h�4���O��/#�;��dR�@�g9&�܁Jh�x�S{�[�^��R��[�&�F�{�I�82�k�XY��͂AV
�>y�@ƕ��h�X��۳*i"~W���rbH�fh9Ё0'-�^��)�vu¦#�I:<4z�i��f%��J���xR0���p�B�X�4���<���qQ�g���1Q
����i����{����[JA�jN��p6���������t���$/E$sr�?��2��K�M=|��k- �u�����u�R�BAkR��	��;�Y��ɝ���2Xu�Ǟ����y�"��Qk�+CʅA��/��K�����V%�4Zi&��L�vje��O�ě�������� ��-yU�_`����R!�nRN�ҙO�^D@N������Pk1/½�ފ*���.Z{�m��V�j5?���ǉ��?4�o\��Kks���n�N�*��P���ƾ�HS�7������S=)�b��`�����}τJ�CRɫϷ>���S��PҀ�&W'$�"F�D����� $f���-]�w�td�V7#.��,g~�*��y,5��s�f�����^�d}��[uJR�^_��w�E��:n�B��g�|wy;Yf��EP%�o������N#L&T�_�
��Y���*{�>+�l�A#� �2��(]�VUwX�aO���!���O���@s��q�+T�{�^��ޞK"��9�{ԍ�{��jN��lCm����9���h(IcY�q�!�W�#5�V�8��Jz�ړ���h�AC2A8�^�o�-��d��;�*�)����.�_n����6�r��kт�45x�CPt���V}�Im}[
/��`R�3}�p�٪I���RgfܖiH�o�i���P���(c}�DNpTj���@��_E��7N51m�M��9�V�O������^f��]���M��v��>2��s�TR!{/o�*��~s��O�%0��R6�#���ٮ~>eX̂w,���Q����� F�!-i#>J��q���G)�M�F�co}��SU��+����KS��L����@��W<�fP���No�]Q|}�&��\���\g[Wjg�������=�>vhUkY��8"��B��B�s���\nO�ɏ+�m�Y�GR��9޷�	�C�������>��`���[P�Q�ž���R�������)Q1b���<l��Gl���ͣR���υ��ZmwK���5�]�?�GI�b�3�3��N���k���0��T���/��7���U�V�ൽ����3;���{�\`^Qx�fA]o��U�qw���K����d*�X��4�\p'���B܊�hg���b%c�^��v
R��~�<L���3��8��Wڠ\3�A�Ϡ#�XROXW)�O�����M�����$���R�=�J�Fj��Kc��ۢ����xX�s(��TA:;��Vq��amYԨ	���JƺN8(Yǂ�l(�%\u�CI�ka���¸#������D���H��紐Ii�G����8,��-�ܧ� �?��_;�z�� iq��^ ��4ό�C �$��� jes�M5���TW�Àz�F�SN3~��!�38���t�$����/7B/��)�ў�(b�k�m�����BWP0ЃJ���n��}�ޠ�ꆐi3ޘ��&�����W�)�D
��cW=b�ն��?߲�۞U;����FKk�vNyd;Ɂ��>���^�Pb|�& �^ڂ�b�ȠvP��]�����=!@�'�Rw��ܶ-�K�m���د�gnm4�t�������
�[_K�~��E�9��-~	�5ҫ��Xh�KJ�=���u8��%D��\��~9��ԵƓ�Z=� �~,V��d�;�� ���|9'���CY��Z��c�ձG=�5��?m���[x�����x����S��7�%��\w���;� �6Oy1���}��p���)����zC$��%jעmQ�)c���%��K�2
�
����n��]ch�~����4X�~$�y1��>@N����;�(���w���=^l�7�7D6�
8T���"��M�N��M��60�$��3ib@���^�  �d{���ԑ[h�}:�D0�ܛ���m���v��a� ��/�6��Ϩ=�*@Z�G�8��+��G�s/y1��?��u��XKh8��o�B{;���R�O�KV8� �k���U�7��y9fm�N�kpA̓�j����gR�H;"Y�n5Q��HHԪ�6TY�t]�:Z-��3eC�Z���`#�;s�ʫ���(Y
���<Z�9ә&���^�>��6�ou�-�_�e�;��J��x�����o&O�ЬE�._��1��jU��.g3��^�U��+cw�ig��J���	FI)z�M��ٲ���%�{&�cb����C��JCTc9�#=��ܜ̏�����rArK Î\�-$]�B�@N����D�A�&��e���7�K�{>k���� ��t*�e~�Nh��,Bny��:���&���T�|�r���O|(�1�����F�.������=v�����7/�azQ�>���i.5��7c�q��9��%O��zk�x��	�GW7�DЄQ��u+e�T��;f&�s�
��?�S3@]Ԟ��?�]�/��=)�2"�����b��*��7<�?�c��(o<��8D#	<"�U*O����b�+��x:���c�F؝_�_y�:�_:Bh�� �hPJ1|
��1��+
>����h��S�:R	zq�X��'��7��g�{��T��H�bT�*�0e���=���l�?;��!忝�V��1&��.$~��t$%�=Ro�L}0B���
stCm,��{� ���&�t�@i�P�7Z���gx�h�>��)��^��6�l�d�Ê��&~� ��Fq�l ��X.���4H���4���8�&���z$.
�G-� ��fGn����-W�?�0#tuԃ�n�-�r�r��¤��IޙZ��v�����>@�`����.�~�gj	ܑ��F��(�s"��`8�����6P�jn��͸�l&7=�W=`��r+�Jd����׹�5�!��쭽�n!�EPK�����^�k�3���Γ���W4l�<\�#5�^���$s��m��i�m�gk0�N"�4/�:!̔�R�/#:�;?iB֫e���w�rh�8P�Qa{g˘oun@��\Z���ݪ����`�?�d���*�Y��d�,�9$h�j(Q2tuY2^��ܧ�ݹGC�P�:J��K��m����U*���m)ɋ�촇���gM VgO�i�ȷ��l(b"���gh"~Ϩ!;+y��uVQ��m(�?j z%]�Zy���\�@g(���6�5/ق��䜦�\,����L�3�<���=��Ռ[�����u�*���2��t�^����h��n�ǈ�R�𣿗�/ﰡ6
�@ض2�Ԥ�Gu��/�c/Px��Я)��N��U��L8�W�ҹJ3X�P��ݍ~&� ��@PF�)�|��rԊ��!�������5�Vc@��q���ZG��t����k��W�,��;�@���Ύ*�?*�b�	i��v"&�2��hW&.�n�P�z��L�f�J�]�;�pL�#ձ0�O���)�uO��^g�-ʯ�z2MP�:��Xѫ�|b������nu���F�ɑ�	=\}Y�Z9���KC���M��ث�t�;�++�q�yr�rz{��L�wi�Y=S��fD3b�؏4���쌯�a�#6��	���o��b�pF �jqhp@z���%�y.���i .�R�cV�����'vB�aO���#���Cǯ�����r���į�#}�u��Ez��x�� W� ��6FV��~����kW�pȚ�mT���G�C)f�d�k�&q����'�Ѡ\�!�v1tc�(�I�S�x(7M4���[t'^3�nj��RQ���"��T��������H#q4F�v�is.�����r�����J���XQ1���c)���L|��^�KA�e-���7�L3��*��j^�~�L��@˜B��R풺#4�bq��桱⮓��@Y��u9Iv>QF�����#����e"�� P����:�L���4ȿ2����WY�2+xG����$��wxe����
eH!��;�l�8���� %�Wra�	y��o����$�_o�R*VVW�H�y"�g&��jsh;V��D��Œ-���(���WTKG{���J˂�r¾��t��A�Ó?L�7�Ȟ���@��}^���}�h��&|j�.!mO61���˓��v�&x�q�_���i�qQ��<��}���+��!+�Qg�뵪��x��5u��Djv�Di����/��\��jo}�j��Kv ���c����	�~����\���J���OZ�?Ge�~�����&��>Ie�ZNV4ƿ
��`e9'jVfؚZ��PUgRv�I������D��j�컱0XH���+ǤϨ������l��'m}�jK��K����@v+��iy]���֣���1l�w�c�m�o�;9��6sQN8kG��.2�F' �(r�\v%J=����9��*�+c�MV��������pr!�}��m�[(u@w�S�:�����rV4W���g�⭌�&^�#`�mA�H���m|�)c�N�D���=<_Ӱ^�u;��O�����S��Wp��}p��/d�_t��$���$��WXԓ�*������`�3�/C��H$�����e����{}�����Ϝ����&NCV����+$0���q�B# F���!��;i�Ƹ����ښK�K��*g��1d �t�?�j>Yܕ�@��~f^ <_��Ɦ���>��nER�{!�S8y�~���)���b�} c�Hx6��?�.��F���p�#�^1�F7R�ۗR�z+��g��b�L�$HF�=���(R�I�\i�e� �6��=�6&��gYG
̵�#�?U��v:S�6|��G��I��^W�q����_c�x+{A|h��/`21�3�n���o�R�Lq�3 ��7_ưe"�d�����u��s�ϧ�-���3��̪�����x�.N�0$�[95��D�눦'Fi���S�֏�[���˥�N�i�����Z������}f�t,n�����Ǿ6��cO��Ց</�np8򪣕>��_�a�ۀ"G�����H>c��ZՏ2Ɇ��8B�����/��Oi�X�ȼm%+J��?zΰ�8+`�AJ"��N5���tp�lz�U��0�[u�A�lY��y����f�Fb�5c����ZR݆g�p4�8���W�҇�\�8�����]G�Z�]0�7��-������FѾ���|��5���U��l2�8̪9���)B�}OcLGf�,�=�}16�$.ާf������7۷�&#MܨJܖ�j2������ҙ{W?�X@�h�f���o�8�G�JdCc9�dH���ʻ}��O��l#�Y,�{����q���9�ł��-xHi�j�:Y���P�����V0���j\kԹ�����]�^�k�B�
E�[��~62���X��(�����lE�b��1-��������M�VQƅ�@HV�N��vٿC������~=��L�Vv[�)NNT��.����ӝA�n�͚���"�����	C<1ۗ0���vח���
=ҏ�	6/��J�:���e�%_%�_Jl��ds��(W�`Ȧ\Ճ�LX@�ũ%kL�B�a�TuP�� ܥg�,&�y�Sw�J��+q3\CY��(��4	\�����_K�$�]@��t��֧�9\0Z츊���lT&a�l��R���&�y]��v>	�)���,'?��+�2�����)� ���X�i�}���Pv�r5�TD��7W� �o�痩����PO��o�z2�"j��.�$J�R.��1��$����r;!1v�o�KbW�§�lC#�'Q��"��xp�P�i��=Mh]�T�&5�.:c��6&�Ĥ�)�xϥR^�.�;���)n��e�u���g��K��IQʶB:-�b�T��W�J�e]���a�g끬f�W>T+5;�pC�'%�Ʌ��Gw B�H�(��8v� �ږ#�Q��S
�eT��)"o\�eF����}��!��Y'5�"���TWg��o�'\=���ղ
�����eIMCm�P)�T�
�'�T���р��+s�/��9ϕh��3.��� Yͨ}���.Nu���#<@�W�"<q0��c�F�F�,��<��0Ƽ9+[qX�CRN��5w���*{����[/�9���2�1�,l���T��~�Ub�o~+�|0����{�l�#�X �k�<+��������}���&�<Q�B�_����78l���(O���E�~�b�O�y����	��G4��T�Z(�ۉ �LZ��L����
.��q���/���X+���'�Ȗz���w��o����sR@ؚ,�΃4+�K��*,��8��g��Y����
�i/+fe`�f��O��~�\O��0;�q�gNؙePa*�i��|���Ӽ�M^P��p�N\��-$S^Pөw."��̠�sϭ��.t��;�L�a�[���/"*4�&Q�a�C�#��%�Rv�x�J�I}&h�g�O�1�^���աjd�'t���͢6�ʿ��떳z���L���D�b�V�+��8�t���ʵ������9�kA����͡��eG�E����:��@]��,�W��9w!*R/�4�wAK1����x�m�&��v��O����L�P�̇��3z���3���D�"��2�X)�_��m����u,3�&~�\�掑'���sH%y��I
��]�5~Y͵�JG7���D�,��ɒ2p?vu�UG�%FCd�Q�*ҷ�u�	�4N*|X|2y���E�c�Sx\u\�<b'ӂVbW^�~G�v�lM�E��C�q`���o7mQQ�ѡ�����X�D��u �����z�UP0d �X��Tn�e�T�ݽ��%��~XJE9_��a�6u��n+a��Go�h&xQ�4ݒ��-��*�A�����,ގ�F@��
I� �x_|&����i�gR����˭������v�n�ƤW[]ƥ�� ^�=q<��u��Å��X�S���`~��6����&���T�=s�����!�QƟ���hU�� ��J�?	O�������,�����s�C}]�u�rP��K�k�s`�^';b2����ݟS��,�[x�>��Z[� /n�����)��uYT����|����+tA-��zJ�w�K��	�RM" ����'>��3uܔ�������@s釨 ������d^ ��4n����SS�(r��&\�汻a��ç��(�Ntb��u�*����	�6u�V��4J?ԷX����������o�_}�1�U)�]90S�I�x����
�D$�m>�-��P��?wR�͙ە�5�3T�K�2����ZBl|1���{�85>����+nx;`����`�2��	w��bB�:C�98uu<��Φ�?2W��� apP_6�E�I��k��~����O��\������FU����k��0Ap3���|��9�l���I��L�������<T,�70�0� _��Q��Jb�ʼ���h�|Q��R��3�Z ��9&�!⬞�}o�m�?�d7�����謷�b��X0L�l -Y�b
q !럝����mIe��������vg1t_��s0��'4�"c;��Cد���I��������}ҲTV�F�V�����,>�"
�����a�d�(��5��B��s����c���W�L�q2q�\��}�8��+gR*!iN�g���󜺍Gη%�
c��i6�~�>��#[���ծc�R�h(�����P��k�M9 ��dӒ�Rn@�bh��m�fj%�]U] �o�ν:�T��`��񃝤'l_bQV%[��Mw�l3iΖ΄���T��G��G>��.�Ȯ��_�R�Ѐh���VU�˗�+й�ˆ�j��>�"gО]_�L!�E����X�P��,׭K�5�M������5c���Wv�. Y2��!BT���D�=�ÀNY�j=��o=M�Z(1��;d�ekpׁNNV�0�Z,��Î�ֶ:+�r���װ=;ޞ��l�!_����(�SG�b�0(A5_�p����roG��D�~���v>��f�M����v,����3���®��c}Q�E���+ԙ�C�(<���x���pYs�-�x#�?�^�7W��A���K�$Up��B�_�2�5*��^`���C��_�K��!.�0�Y�����3���Y�:q|�蛭������t�OZ��l������:A#�̔KZ�;��3VD2�l]�Xd�{������E���VUC�IpRt�4#�>�mĝ[�b�T;^�>\}�_���
�$G��#��;�t[�"�W�.@�\+�u}�|��&,s1|�U�|뇱�Ż�#�o��jg�#D ή2m��;K�6�
�����;ƍ~CМ��7��:-� 
24~��Z4!48
ʁlW�eJo��S4�YfX��*20��4�pF�.L� -n��<֧܄p8�eל������qh@b����8�K��1�1�z���P��l�z��~�H �DNN�ݵQM��d�COT��f�#�9��u&e�~��zXH3\��1G���\>�@k�R�:���Z#��>c��&��������B��L0�>��8�\���f���Ӧꯚ��OT4Qg�0�h^������&��p��x2�Üh6ᑓ� Q@��w0[,&�[o�?G��N7N5TgϙWk�ĺ�Q[2�eCw�*���U��:��w&��
�>1]�� ڦ�q�#]�>�ר����6Twg��,�U�9W0%[:)�b����2�����4�}l��xj}��Nq����i��n���@"m�K�zA�ѧ�NlYQĲ�P��R��(�5�Ȏp�����d�����p��1CDA��0����X|"�9��cE���0P���E�c�1 >����lTa�w���@�#Y�߷�b����n��Ȥů��ǫ����h�v�±[�zK4���`�<�����^y�1�"�	���{��FL,���tT��'��������H��8��ac���\�)�璕�v�Y@=��q	��iHSؙL8�p����՗��v:I���o�lV)�K���X�]?Hг�	=��J��NN�I5���i�k6��:5Vi��ü�4�h��O<�n�xC=�_)vs��d�U�A,��;��s�����]�>*��:`s�3az��%��%,4�qs(��N��~/�&"��>b�ѐ���4��b���	 RB���<�л�L@$�oIO=���|I�5촊�3>@�4�A;W��f����T���x�
,$�����vQ�P^��5F8���s��
i��zmN�0�*�E����Aq�5�r����!\-�~�FI����P~|��6^�/�BU�g��s���{�
 Ȯf0��)��W��b��4˖f|y����%Ă{+�naMQ����s��x�Utћ�5�w����ұU<�LSCλ�Z�ۢ�a��G�� 0�̶� $ɖ�%�8��˭�Q���~�+m�Y�{���EA�J��0��_q,���#�������V6��N*��=x��{2��GD|]As�i��_�;,VU
	����=�B煳�Xy�j�Qs��H��p�g%$��ꮒ�Q~��MpDI��3閃L�`�dj���,���֐0K��[K,=�%%?N*����]�v�敖��;/��T�-��ےR�]�������"g�;�D<�z03���m��	��q��I���1���WV�c*�w_� s�޷�Ez�cA�ͧ����h�����hB)����6G�5lH�j.�]1�iP�h���7WL����M�M��#�ȏ/,���	��+�B�:Ћ\�Ռl�-o���}V孻+�cKF�I�k�e�X�S�-�d`�	�°C�|�|�˓ӟC�K	�|�"���3Dm~Z�L������B�� ����؃�����8���|��r�\�V�YH�t����by��3�s�0V��~p��u��1�'��:���1���Mt{�W~�&�z����	�[�_8B�8��o�� =i�n �-{�a��љ]e�ަ�2�g����z�-�T�����D�����W0s�wT�鰘�J]��*}����%�ʁ	��ޗ���_'�l�'۷��gb	W�^�[��c%����w�%��?S����+�%��C\O���ܫ�@���m'ob/H2v�܇�M�kc}>���l�q�L�f�S�e�̠)B��?�V$�4��T��_t=�ô�� *bA�-���xN����b�;�-w*�y�ك��b��̠�o��R@���C*.s�P�BYC��W��=�)��,"�;t����Fχ+�u�>6�w*���¼(��nN
	��5kY�A��n�����M�h�K�]����=۽��V42Aiۇ��!143���������� ��CP��HWDn6�Q�c�$����C	���[Q����{/��4��qOyI�X����F%]�n���L���L	�B�8�I��̀��:���r6�Ȋ��)�_^�k�|c��"����)6y�R5��q���װ�_�^5�=�����YW���j���5d��#�؃}_�ȁU읤B�����C7�j�;e���� �miF�#qb��H]a}�D��#ܑ?o���\�G�>�>����v�C�x��/
S˛�����L9n�=D��*�u�[��j��s\���bR����Ę�l�l���J8�v|eIΈivR�}�[1�
���E�d��3E�k�2��K0z*H�&eF�D�T1ޚ&��1���k��=5g�>`�ݐ�޷wk(�LL���������'�0���Ȫ�$�pz�	!��ѕ�$o� ~i!3�q�>���Uʥ�tV([N�*y�"���0�AkR�l�q�GS����u����d;N�Y�!>��5_�h��������*ViE��\�!=���rd�	�E��>\��!���??:�)��GXj)t��R�mDTTS]��Q!H^E���D����w8��������Idރ�'#Ud$�/O�6M�����ˮc����N?���e|�O�u�s�'�A����X^��V3er��lNy�2%����n񃫫d����w �q&C�F�ҵ��,�����I��6\6�*k���MG�ƵY�ƒ��5Z��#"�!�?���f�ё�3[X��|J:��2�7�ch2��		�UC�E8�D+c� 7��&��=�+j�0� UR������O�VT�;
��3bTU��3	c�5a��[�I�`�y�����Bl�^o�=�O�JI(��̡��18~��ڱ����Gk#���R!�Y�D�N�Yj3�'����0�f��1�M����D4�P�X6�C��7	`O�ܘKՠFp�G�HQ�1ǳY[���;���� >�?�Aq�,Z�Bʪr�v�趫����l֌���g���d��=ǐ�f�Ū��!\y�]n~CY�(�U�P|�R����`e��V0��d^>U�eE{h�c�%gV&���a񪥊�r�(W��z��ž�k)��Zgp���Wn�ӵ�ݎ�D��f� �x���e����`�h\�6GP(d�E'�zv� 9Gz7����f'�i��� �caϥ��S�ͼ�����u=3��u��'!Q�ڡ�u����E�����`�=�O��|�k_�ƃ����wכN����g���C��.��ެ��zwh���q�S�HH�Z`V�U*n���72�/^{�O<|>�C��Zr�3	�v3ZG3�;�L�� av+���!7Vwj�
h� ����	4Z������P�T�gV `{|��O�)i�z�2���F�j�Dcҳf�OJ�9�`��M>r��>/���R����M�6�U=d�t�!7�==x�IT�9��5��ĩ�IdI�%���*&X�_?o��
�"Ӹ~��@S�Y3��U׸���/:Ul�B�$�PLwc��A���5�K��Ez=U�̄J�����������զDn里k�-���*K��W��i▍�1���2]:t�W�6^ޡ�P��O@�O4,��\ �s@�Z�4�/Z���5�g`%�c,�E�SxH:��I*��v,D��ۗKR��$��$�;b�K2c���Y�C�h=�uKʁ�?��t��������M2�«��%�Se%�߃Y�������&�W�3����↸>�(6':t4@	�r�o���+�D0
�0"A��nؙpa�;6� �^,��=���A��uwZ[��Dd���h`�m�iΓbWGqc�4#�9�>v�=���Ai�$Y�a�~�)�`-�/����^߰�wW���y�e�����j{W�
�~���r��Q�k�2��;�%ޞ�B�ՖJ���#�j�VD���ssH ��=Kq�+�m��ۥ��>l�Y+��qo�~^%��鸛�.�YԄ�1fC;�t>LC5⌁��1~vq��B��F@�7�
Bª���߅9p<NV��%k1Yy�;�HHR2�Mx#�0zF<�qAih\�>�j|��]2O��1��"�L���>�ǻY_E���Td���v��'�U�o6r��9�V��h�!P�&#���$ar�Կ�^��70bׅ��j���d��9�!���dmz�#M��� �ц���aO����Q�+�MOF�Н6h6��G
c�g5Vp�-��K`��9�������հhW��l'<t�a%�)r���E�]�\���_�����t&8i��t����C���!-�Ǥێ%� ��?����(������swm&�
�i�va=G$�/ec�͸zg�c����o�9��>����xJEQx3��g&d�RL��E➃Ưq/L���R�����A�GR
�)V��G8��40�S�f�%��ό����I�[���N/X��`&��|��TH�q�@̊-e#s%�C8����@3��I	r���#K?�F��6�#��xw�5�B��-gF딎'�����[J+�(_�?<�Ă���.�%��z��=�	��r�vh�_x|_Ǵw��b�36?��j�����P�c�y9�*�Ёr� W?�LI�W���	����%K��;��p�R�V:�7EK�ƙ���)B��Y�Y2��Pc��²����Y9N5|&��¹�)5��ե<�8":4޴+r�¹��y$7̙K�+Z56M,߽J�0�V��=�ҙ��C��p��N��Q���[�bo7��]�Jm��ԙ�y�d�N{�K�Sy�L��>(��������-���l=��N�\�N��Ď��{�T�.�K���]�g+��Oq�I��Dd�j����N2����~YZ�>J�eo�/���Ag�^溏-@�z���(-��xx@& 8��X�	Lp��s'R<��N]JL`�Q��06�*���jb� tו��N�
�h�[h$�[���m��C����US��2���o��n���J������,�+���Q��pXh�rSi��Od��#�Qo���{_��m�@#l?���5�7|��q�Dr0�i[k�z�k0i�IavI6(�4�΄�h+��EJ Sӳ`����:7X!�"g�>��߿��E�[$�K(��ѧ�n��1z�Q�0��o��ܲ�F�{�ϼ`Ҍ�AN�sE���j�󃗌w�M9��}�����ј�J��캒)�,��4�f��`g!^hʠ|߃z2A������Ka蓥��L��!R��t�6y�����8`���[�o���(��+�;� p�m����g�)��ݙ�K|#����f�?!F�7��F��������_��,"b2���.�&S��ߡ�O�ٻ�P���͕��4�k�#B�p0���]r@���#�_�a͡�վ�����d�Ǯ�2WI�q�|��Ub��fX�U)Rx,��5�}�)��ຖ����B�2�F\��Gp��a�����|�M /	^g�I�e`v��\�
x)Ǧr4�:Z�"��oz�g}��)����2vj}�c\6E��/��kk{TȘ�.�<s#m���9��h<�ɑۈ�n_�iBjs�ܮ�s�AB�t�|��B�j("�����\�!���A��q�%Xw~�JU��>1���×�nk�vS��>ԨS�Vj�H�˿N�z̬UC��jv�]�'�|�(�b|�F�rW:�����*?K��q�M������_���^Y�cjVy.g��`d{�ɜ���S�NjV�����L՚z����~Y��k��n}*l�޿Bk��]%�l���׼�2\>�*���G�x1��;`��d�1��k�#��K�A���+���<k�g}��}x*�� ����I���"ll�\�r������VҰ7ot#���~r���fD�>m�
��`���F �X �'f�2ٷ�X@� q�#�&
�|���9�]�)>�ӯc^1d
��/�r��6{~�R��)˴��7�,R&:�������5���zt!�(q���vX	gz��,�P=MwJ�@��,�������������)䫈��ɛ���m�$�@�`�I�����]�y�^�t�>Z�㨭{W���s���)�1��܌Ԙ��H=ve��b:�ʊ�z��ѐVuu��%\�HS$.�r�.�=2P[B�f�e����\4�0FLo�?�S������%X8�B����!��2+�</�~\ ߼!�_�u�am�_b{��?]`H!��E�;��KI�S}w�T�i�N�8�A��8�8�Ҙ��[�~-�0#2+v#I\�ڮB��<_���3�b����j�DNnJM�h�ee �=��ş���3Ny�r���� ߺ��W[��c8\Qًe�=��G�,I\����g|��O�gF�t)�N�s�:�##4�BԷ�p<��`�qD>�.,:��������<
J"/�\�"��a~GӞ�?|���� ���Rpb|U�;2�iBb����.݇_�(�o��cL�~���R-��[��	ٹ��u:c�7�$�i�&����VD>�������jq7̒YF�8���4&^�K�&�fr���v�qH4i���O>��v����5-���0z�n�_�	�äÆdk�c�#T�G*����.������U���<�\��)��}i� �g��p�{ �^:zZZPE"�`�G(�f+/.�q��~��Jd%x���b�7Vc�Y����n�=rzvu�M����-�O��'��ǵ$i�N�������RP�����֍��̈́�s<����u��~<�J�6�묫�C"n;�2i��z�4~IҢ:��Ŏ�z��PcԿ�Ȱ1
�����Վ�0�ޟ���A�E��q.K2��ü?t�b���0\]L@2�W� e �o�ʎ}Y�hT�b[��Abt��u0�.��E��UQ+����{��j4�b�)��=7��~ع����H@8��u�9�,7)�h�拤/�� ��鬤�(1y��jx�f��ZRi��CN8b-��L\�x�K����ƃ~�`�Op�!���<%�p0K�\�ԙ4�\��q�θQ��6��/G����g�N�>{"��~�h�N��5댁O?�5ξ�K����}��j�o(EزC�5�r�m&��Ŷ��M�n�����˳	��n-	s�~����sZH�N�J���?���P�N��ڗ�u$����?ˀ>���=��c�R�(Lv���O+̿T��y�� ���?7�����JAm�6�&�ASN�/�\A�{����U�>z����JI��et����i&=���55&�֥4���wj|���R�a�_R��Ƣk�kYӔ�����j�Rqh�B�V�+X��4�mؾ�A�Q��jϗ���1��5�d�����B��9�@i�� ���chIk��������4�]4�`��!v
�%o[�	�`!�DD����?��(n�[�6�\�hW��r�5[v䦲�2J|d��R�DŁ�t(WWZL�X�.R�W��/}s��M���,�l?p�Bm��E ����@�_�_>k��$�\4�~�!|���~Ո���eKr�[�t0��|�U���ԣ�����9���	�|o��z&9���'�-&a����V�T��kI�҈�<5c�����Qt����2���kH$.���xQ"���39�KVTW)� ��^����Mؤ�X�ɍ2i��녍L���HƜI�LԼ�j��F�3�2%�A?��[P-�<i�|I��a�x��d@z{n�ut�X�X1�����I-���Sܢ�J9,�Ԅ��[Hk����As�R_ވ!s��]����יMS��<��t����G>K��L�4���4^te>0���E-:�!d��{�[�*�z&����l�w�{��
�[A�&䪆J[��Y�2EX�Ŕ�4 h�9��F�9V3��i�X9-F�j�8�K��l �DlB.�R��k�e��~�!�<��^ۛ��O`��]W��Y��Z?��A��!���||���SMcX�6��] r�����t6a����O�3�ח���Wn�,OЬC�.��XoL�]R�խ!�#�S���l���t>��/_��0�pN����T�i1j�_��!n���YύS
f:�x��I�*4��S�lqgW�)�ZW��ר�a�O3v���i*����{s��R��g"v�ۣ׋�c�&�5um�2xNT�[12��JHId'>q��C��U'藌l'�I��}������$٘/��,j��'�L��!瞧���O��H�ׂ�D2��r��h)"���Q�L�;_��]�nU�������us���}�5cӲ�Qbh�=�4��M��K��5�.��^����+�G>h�{=G�QÌ%d���<�Cu��� c㼙��_X!�emZ���7t��^Rt��؏֢U���C>`lL�_���׸�
}�W��Yh�aO�U��v]�@�dj,����)!��2QQ�1�c1�)-�?f�6˂jQV���S>�^Ry-I��$��%�JU9`a�Ӣ�΄9��.��8��m	D�szlԸ\�`I�� ��o�[lڻ/F4�JW�w�H/hA�=MUNl�P�s���r��m�m�z%�U�"�m(M*������S�dg
pܔH���u�I�=�"���xˑI�%w�2� 8E��_�KC�*�â�RfR��Kɶ��Y�yF=���=� ,l��;nA��}���)^�u��Dg8SՕ({-�A��tm�2Yp�l�<�# d(^D!���L?���rR��8��;υ�U�q���k$�S!A� �H�:&�����K���>ҟ�Y.�J�����!d��;��������:p��3�d�� �.���y>~��T���9����}=��Dxy��<PX�����ҥN�5����c�wT;V��ܔuO}f�7���	�T��J�ŝ.���~*�60���8p������;�s�^�`1��P?oQ��|H�z�=�%�4,��Rc��f�
?��],�BWτ֮���DJ�<��g6b����ťٶ�Lu&��·�.X7q�;cW���s�f��ٝb�]|&j�ZS���x��W���G��71���۶W�3�˅fI�_ {���;�O�������a i�e_�	�(��ݍ���d|��5<�jD2=c��y�g�����X���j�yE��=����82x��k��60�1徴��~��)�$��V��_�����I�J<�"C5�Y��M�̣�oO�'�K�P�w�ݛ�#|E��hCZm:\TW�o�X���j��É׺�+�H�BU��
��;��~^n��!gOH��̃JL�5)I�;ߙ�}�j̀1�C��P�C���b{+9��ad_F�{��a8�5/��I���Y�"�O#T.�hM��?�e�ǌ���X���%}��K�C���N �uG����K�#�\D��dʻtÁ�	���� ge�M�*��c&��<h̹�Ce>����7�^G�b�b�)�K]�pj�?�K�6l�n�k��T�ޛ8���eR�����@��_f�L6!�4W�)��u����}r��UO|�gL��X7�����v�ٯբu��V�b��`r�?V�=/�m�GW�s���S�&�j����bB�H���=�v�R�� �7�N=~�2I������}�B�S#h2���p�Ŵ�O��dZ+jf�ה^ 	V��ݬ�����KӦ�\�>���̈́�U�~l��灂ɋ�C���8pș��WE0W'�4�6�[26<	kY��6&���u1��� ��BͶ��#�L]::a��jfp��Yj�+�S��m:j���� 3��Φ��ˊ��FD�bU���{�-�$�ģt��	&<�\�ٔ���B+�^�}���?���_��t,m�U�����>�ec��gd\\5]�)dm>�0��w26����N�Ja&��)0������`aq���eͥ��|M��{�gR-"�Q>��в�����e��g�����	����9܍#���t�s�m��=Ɗ�2� }U�6��i�]�9�Lo��r(� �`�Ss���R訠�:sx�/��G��I����e������ ٳVA�";���d�"�IS&9��%�y��Ef>a~0�|��f�=�tL�_������WI�'�� .H�>��n�b���ѩ�M1�Z��T�/F^�f�Og�Op�NJܶN~P��F�hI9�_���}�s��Y���������s���Ϲ� a���H�R�_$�8�� ����5K����D&
���;CPj��Ǒ� �e��Hv�cP�k���ѱ�Wx7֨!VPL�]�n�yh�e�� �@���5ú����=�t8J�ȯ���e6���8ܻ	�ũ��t�=����4�A�l�cql�Ԍ�f���b����e�����-5�dΑ��r�t�PX�s@��# � �@!��Z�u�
J��HP��j�&)X�9����Ho4R�bVWc�� ���m��_ⴓ�>(�E�^�m�ЭnR}�i�;RBaM8],V�~!��ڜ��e��@�<Y�(��>;��rJ��K9��y���<-��m�C���x��)-#���0���NH��P��hm3��y0\�(F:�7#sc�ACY��?i��Iy)X�CP%��i	�D���L]C-S���q�mQ��#̹.�EC[VW�__�!�6s�t&[�E)�?�������L/�����G���AG����u���2ٰ�É\��>\�����^S��MMɥ;�� �����#u@�u�^x��oG7 4���,�4���|���73����.��G���bH�A�M�W��I_��Zze^VT~������ʊ�H/B��7g�x��fE��А�������۳N�P��Y}��֊��ZȞ�3�2�0���[o��E�z��؅�P���
�V���x>���J~���+�u$�RO��:������£�)���q�(��T?�����n�"x�0��@����\�:`��+}u0c헷�T�FT*�#�v��*L:Se.�F&,�޾�_�'��m�E,j�'�=�����J��C>�Q�a#2V�۟,�)��|�B�Z�tc=P+(����|���_%�DO�M�D���J-���9��|���\?��B.+��a�yZ�?�;���N�|�J��!�KF� D����|�]V+��hM�/ZO1���a��&�e#�2��vS�q�d���φ��󦷰�O��9�ۖ,�}s�׷�)�+i<}.au���k��ۭ�M�K��Ry�*}5Y�c�׎UB#�m6����	����UX�1.Xqˮ��ZW��
��<[:ۜ�+�5���L��C�!��gb0�����:L�� �(#�4�x�w+�m����_,N��Q��� ��<��$�1��Ej��=��/��>l58��Z��e)��=`p�+V��o�����T��(2kP�4~"���f�&���P�_Rk �%LBH�bYf���z*�=��@�PFH���&|d6R���%ݒ�g:V	��$�Ǘ1�tҿ����+xS�&鎆h�	Φ|��7�O<9nМ"��k��YK0�&%��1�̂��ھ��ݭܢ�Ejy��|�uV�g�1	���.����V��{�2�qW˂/��T�YP]��J����]{��><�_y��|��z���?��%����81��Y}�w�w�1G8nY_�)�a�S.b�ë{��)J�j�N �K��&A�;����J�[��e?�����z���{�iM&k�z'.6���x.���m��������W;�9U�@o��r���{�
w,o��"����[
{2�s�<�tK=/ƒ��
K/� d^���[��	y}�#�m�)]w���JF�$�~��"&�v蘆-GQ�����I�M*ߝBǒ�n��|��M�p�n���O��D!��j�?�����3a����(� ��ӈ��	̪]���)Rq)��WծA"%rnM�c��~��y���S�LQ���R_Yzb�^+֤°@P�d��@����#�3��6�1qk��&�ؼ���;4���<�����+��6H��Ứ�ڟko� !X�T`B���CB��ؼ�&�zM-��4�;�I��߾|7
���ܳ7�Vh�����aB
�{����%Dg貖��Q��!��mm�����''Z�ӓ��V�)a9P��:^�Z�����_�y�-�}��\�Pc��²v�Hѽ�dX1Z�����1Y�Ƚ�؀�_�R�i�6���u^G.n2�v������~�AG���
D���Z�9N��=F�CX`�� ���4Z_%!�SuW�-]�n�I��1�B��YMC�H��~��`��נl����|\M Cc!d�����Jj3#���G�KT�ÒоN�3C�0}Ii(�M��ݻ&���ʰO����φ8d;�(�q٫����s�Z���Q����\�s� �8��{6I4H�����~�.Y�a�����kЛ�U���p�!ˎ�|,Ω]6��1)���p-��ȼ0����=:"��A�ݣ\'�8G=6��SE{$�� �1=���jX����'2n�	�_�d9j)��S$`:<����_���5d:W2O�a�팾��G�~������7��k�(ʦ&���7�r�`�ʌ��Z�
*���]FyO�u���q�zuk�L|Y��ֵ�[�-��1�ys-�G��"Z���[���Z0}��Y)�0������Ħ
6`H��S�D�]=��\�l�j��_���m���mE�&�I���Vr�L_e�����/ �{g�������8�O{>1 ��z2�a_Vl���U� #�(]�x�V�:�����dÐ��p�du�4�[�����^����A�,�!� ���D-=�QF3v��ݎ�~�Z6F�ؼ�p'�R����������>+�� F��&�� �cCT����&B��,�i3������w��V�(���J�z8��oWIxc3p��>��n c��$����*���=p7�K@����Ď��,�@`�<��x���{'�� ��n�E��s����<�r��֡e�xb�6��z��-�ph_���5!���n��v_SO�,�c�h��k���� ��/��ҕm���;�b���.��1�U�L{�pV�ߋ��rr/�;�T�Ea��cB`K�_�;���lןV��O)�S?�(�|�ў�S)�+2�*2�I�i#ز�8z#�Nڿ����_�{	8,�D6�	kTY��sd� _2G��*]������)�I��m;��� �6�'�
$���~��D�c!T�\cB�^F�~'z�G��l^�i\�q�;�->{ԝ�i�4#�"��>n`8��&G�8�v�u�9?����^��z�_��
�Wy�+>�JOuk�JaJ��9�>�⽢Z>�o/\��Պ�R��~}�I�#�"?�k�u���fb=�����\MƯ�G3�9��HM%��f����/<�����f�:&��"{H�N��A3D�jCU�V�xW���]���� 
���wΜ'�}���f�����Ԋ��Џ!-/���*��m����s��A�i�"�l~K�d*:����ܦ����/@�����P��p.�C��[|�Q�K�X�
�s�{�e��k�w}|��7��-�O��]�D��M�w�.�*A@gc��4P؜�BZ�w�e���Vi�)�<ܛ��k&��;Ըw��Ͼ&4��o�-d��EHϪ���
@xa�VFؕ�t�8=�Q����d�Tc'̓L��J_6�_��F2d�R��K��BBٽ&N�3���:�&F��s�vfB�\p���
�����:��H���
���8N�i��W������ x�����R#��	9��oF���nۄ�v��~|��{~�ft状�}Vgq3�oW��>����kMz��Jd�H,D��R�<8;�Ѹ�>��A7��$�2#�#��|<F�>p��]�8(�)S��q��$��q*��7�䣝3��(�Ҵg��tf��?I�o_���g�"�W `��;�Eˍ�4�i��Hb���_�n��E1����O��I6��( �
���T��	ר�WG�i�Z�=^�a,r0йM��p�2}N�}����
�w��Lf�*�aJ&�xw�������T��⃩��jR���w��`,�:�,�}����U����4N��.`���h�G�Xj����WC��$d�(��B�WΒ�6�����%L)�R�A�\C��x��+ruC	Q:���s�*[ʙ$ɲ�:T���'����,�x�ҝ�Hf�Tp�c+��� Y0�N�k9u����@�\��C�a2@*� ��ZUp�ۊ.�<՞�`P��6�ʽ���������)0
�b3��TN�a��g�{ÎaG1��9t뻳pu��Tʉ�uR����A%��^�}K`7;���Q4�v��E'�k���:;O��y�M��9
p�.J��˓dz�������Ěq�� .c�6�� ��7�|�X��'�J�?�v"��80��Ѝ�h�3�z�nS�N��ȏ���	��>�6g#l$��4F�a2F�!ݐk2�Gs
�Lr�����Y�'�e��U���C��l�A�M')9G)8���{�V��Ϥ�g�����-���A~�8{��i���ul�1�|ۣ�	��] 3#"�
�;a���փ��2HUJ�nͼ����A3h!	�c5�԰}WNs���]7���!�V�[ͧ�)��b��`'|���+����_�M�U`'5@ �v�Qpώe������$~8}V�y��`���{�a�ⷝ�g�� :�k�U��Ӳ8��jI�݀rY�p�^&�/$/ĳ���p*��	(�����O+��|FlV��	e�OMG��F~��p4��2�;��&�5��}�����N��5�l�8P�#�QB=\R�%� �e�m(R���RR��b�S�9��g�O�Fte������1���J>`�V?���ö��Ī�<�c����K	{�L���jO����&+��ϕ�O�����pe��"��K9֋p��&�=���� �:���5�&3ئ����	��W�����%���I�DS�C�$Fx���C��
���O�s[�կv*����`LNh�5��;s��-FD*�c���Խ5����<�Jc���
Z����9~�c�H�[Z�G8Dhw(�0s'����M
�O������Bg�~����/͡�M:��:+O�Kr��_E-~g8��,7�\m�a��y*�v����$����Y;��V]!��/�?�5��i�Ñt�a��@�jϘ�ro�:�Gy��)�`��d�@?N�ڏ�&y��l]}/f/��q�����ޫP ,�bID��F�x���n��}D���q�T�S	����&�ڼʹ�q�^ȕ���5tl;��X����e�T~���!���5�ӟ
�V�}�Z��Gw���^^i��"ͬ���J��"�ّ�*�V1`v���cSӷJ�-%��Hr���W���ql�{HO�Tگm"�D^cM�U5�4�f�+��{�@p�{y�d�!
�)=����S�m<Rc��.uRF���O4���<=�����s=_�UF}	�u:j�8���C
��1��u�kU��s���I����"�*�G|�IT�a؂�9>w��qx�|v� 	)�Ƃ2O9(走~�ma��XT(f��u�'����p�Us��;����]�@)�����k���^Xg�&o��&d���p�Vk	��@]L�DvX�7G���`�/�Mu5_�'�����'3N�����1��v>�֟$e]��I��'�jͣ��)��I;��a�`��|I2�>A�d��aJP�\@<���޶��\��89�o5d�^!	���E�:�Qp��U�_=0�M'��IM�ݬ�lݴ�:���ɑ��?F�IQ��,J&@�Y�|�t�<���>�$ �
x`�<fLuG �ǯ������`L�[r<sdx��� ��w-I�Mx���e�&G.���_�f�oK�nH]s�fk|)@�q�`j5�%�H�}rsQX��[+�ES5�Y���"*Щ �C���٤3;����o���-D&"�X��1���`Ñ� ���@)(C<�"R�$���/d�S�&4�V�D#�K�����l�[�ʊu�����ЕԔ�^��պME�W�f�%��I8��4V���Kb*����Li��bzr*for�Є��b=��Ӓ���O(b]C^�:v�ݺ[�C:�5+��H�RB>�$��2y��I��?/<�.� ��8�$��I9�fȯ��0��O�yS�a�K�Ԗ"ͫ�9y��C�+��ޫp�������������׫�-�6�`�>�)�_�I�J%���ZӦ���'��x�n*�LT����\ӆ�;cc�Dq���TF��I��Kt�rluܮ�b�����M�J��&>��-�H�8��c3��uي`�y�(�$v4d$��u�����z��zG�#%E�y-e������̞H��sA����+���w�G��[2�����cCk{"�Л��$���^��T5��5#:���cp�؉�>��))B*b��0� UF�T����,x��!�`�ry�dEC���|�D����L�������P�2-z=8���)j���z�(j�#|	�z�i�y~ՙ���chL�k襤i�y�_���h�.���Y��|����͏Y8��L_��jGw������������d&cp�k�!��I���lL\fh#��t�>�?!h	��u��t�B��q`�(>��Vۜ�x`��ݹ%��;�v�����m~�D�l;�uK�D`��
�ts:����!sNoE�W+�:.�a���\;�w�B7~�k���x��|�4��� !�4��}[a�ؼu{p7��ק�8���B�p~�UሰʝB[�`��(�5���o�l�&|!���$΢�G�c�~���C�eT'��5�cB|[���24��\ԝ��h �T��d�$��4�٫������k=mq�-�~k2�/�zn���J��o��[�KNx<�y;�%���M�AP�����m�o ,��\�15kF��K��o��e#k�G��3E�+�M�gx��r�f׍�AqP�v~\ 1fr�10����ʣB ݇�m+hz��Aa��7��rr���ؑrĵ2�1($0u�]
�~��AVZM����w�f�b�D
�\��س��#GVwl�VLk�$ґ��"�dÉDb+2������~cp�!����p���/`��Z]/�N��o��mC6��3�~G� �@v.��r�"E� H��Bz�u��W�y%G�}|tXv_/�=��1[����ܪ��w��q~��_h���9�&�ū-��&��� %�	�΂7C���'��@x,��ax�;l7��KdL���/�����*^`c������9u��$�o���1$��l���tn��^�D�u� Y����9��$�D;��"�r�.�Fz�v(�]2�@�j���0-�.�]j�����|)cե<�o��q��C��ɽ�ӴʥrH�mn?��8��ؑ��8�^�{��%z��.��&�xvJ�5`�����j
x5�Ĺi�������eF��R�a%.��'���=:V"I
jX�y��kJ�>GO�O}��\��,8��=��Xw4LQ
�{�:��ϩ�H ��?���+f|��t���>(Z��u����W7[���x���M���h�آ�^	?꟎hLݵ�4�,;�=�E�<�G�\�mA]m"�o�]j�_h���UK�i���^W8��'���$T�g�c~��������O9ղ�x���	B�Ȓ�X��Iڸ�(p����uO�|X��Z�x�G�M TR�j������sn�<�\�\�O��P*?��#�"a�ރ,�$Ė�Jܹ�Zߓ,�"�����}��ֳ���YL��$��u�x~��	-
�l ��R��h�i��w�V�����x���wZJe�rYv�&��)��@$KJ�\����i��Z�(�P�GD���B�\�1�L��>�.��#-�"x������]�	)���"N���V���Es����2��6\i�\a$�n�P�'�z�_z��	q(�(����!�[���N�����L��J�DT-�B��f�c�e�eC/�0�FH<Y4���#V���C��'��1�9��8�VG��eֽ�
�4�F6��& V�ğ1�V�R�؟���wB�p*���N�CW�S���y'�iQa�p��j5��|����|(_}�x�yp���#T�yI����|�U��P��̓��	��"�IĄq�ƞ"t!sڐ� �gD�ш�0wd�jy1����@ſ	(�eOk&:0�SEA<��e�<���a���)o�4�n��#p�$1�6WR�ׂK�D�Cb�-K�[�
��Z�7s��%� O�ǻ̄�`�s�7]�>{�H�՞3�kuR����<�ScT��`��e��<� ��S,�n�WOg��3�<q��e�0G�/�H^5��Ü�1�K{�
�#%�v�to2���}�_T9�C.�o#�Jc:����ȅ�/,�|�C���	G!���~z����%�iľ�bT�V�(B��bW�t��Ũr��/ߩ���|dwO,T�9�z���ls�M����]��Z��n�� =��T��v��:|���J_^Zb�*A���y,�bn�z�bf-'i�od�'�'��p=��%߃-1�����6f�jT�Rҡi��6�+Ϋ�~�T��oH�-P�x�>	ӵ�6)�gi��f�U��WL�4O��O%��$�[��1���H�5l�Ә�-X�Aq�⚿�V�UΆ���&����j����jD�x�D����.��'�%<WH0S�zD%��)ht(�0���8��3�9�q�CT®��t]������X{�sDY"��[uN4�{_���]���
i� U�'�;����K*<��'=�}CH@
=|,���|X�{��9��$h�Ή�Gz�H��{��w�C�!�?~N��i�ec�rn2~���t�y���X���fX��m��h\c�wz�X�]��"�h
э�����VQE	�JJR�eʞ!�bʱ�j�̀���2��������C����M�����L�n��ʠw�g,�W?�%όmcz��#+İ@p�c�j}?����BP��pNukd�Y���TDށ8����G�!{����N�:��	OM�=��ژ'v�f�W3����<d��IZ=�y�ل��yV�h�تfՏ�nH�����^N�{3�p/(����~�$��5��fv��0{����9K�V�/d�e�`��'�3S�I`@�ׄn����u}�^���X*D.1�p�Bǻ�����vP@��\��?ab6�~Bj�"�7'���C�`1Q���x�)�����O�҇w�rie��<�F��h��l�0/�o7P-#�T U筭�(z�#�@�&��!�dN�1��*h`�6�13��o�9W��1e��H���}�f{qV���:�gZ-t{-g%QC;�2P�l�[q�Kqtj쬯0*���a4<�������%��Y�?8�9�r�*zӯN?�ɣ,����b?!?���%�t1�U>�ӻl����x՝y���DE��o���`D�}6J7�C�l������?�2(�r���9�߯�(�0��}d��S1���+��A3hW.���M�'�R����L-w�lp�\`pm/�yTa�Q$���}1��4�a���:�C2(>�4�l�.q�z��Z_�Ŋ�$���!z�3e=�����(��r��3_7�O��l;?����e�-�_E���B��U�) #1T�ذ�M��&];o�vL6($e���A�k~1X�3!D���<t;n�_UT�{�R�h�H�\53a�'�(��i�=#��d�W���~��;��{�
'�.����d����~���~�=��|��()�a Յ�����(��:���)����9yE]���k���ȣxFH  ����ɜ�N\�}�빞	{�����E�e�/��V
�P�	IcTn{� �t�SS�0�V��{*���K�*�=����D
	'OGe�+���1 %���u���c��e]v��gE����d-D���(y�����0��!8���F^U����C�=P���k'��Z�Z�<ԣ��f �u��mI
Е��F��vc=%�� ����}?�^�#;-��O��ؙ�ݺ��0IކX���;���q��f�}���������j4�r���l�(C��/���.+�1%�6x��s�( ��{C65e`�J���H9�PK�pB��i}��1�窋�VȔ��H��I-��0���_����]]8��Ѱt��:$�Ĕ�s�bv0��LyК ����l�!����R������I�_����2�VF튎����a��ЬH���'����=N=-�"�Ο#���a-Ü<» G�8NQt���+��@8"�|�օ\��1fG�c.���=�l����GE�+]p>(���3��A�>/,���3]�!N+n�T@�^�~3Qt87Έ���}_�.�ɕq���UY�����f���������$�:yzs�ZKvOp�+v��ۙ�I�Q��v��A�v��~-����7$�и��t�S��I�n鸎~�@�'��җ_˚I��J c�}��SfͱR��] �#���T����W��N�JL4J�(t���j̵A�9���^�	�NY���!Y��sBg�r)�v�&P��S�ȡi��=�^^�,��������v��w�i��c�;xƊ>s(m�A�q�Wg�>7{x�)�v�jrQq7]�]�Gy�]���)�;�eY4��q��JI�VH�%8z^J7L�����q�ʌ�ݡ\�K����,#��5�8����o!f�w�d>-�ĐCo�ju��X-dR/*���L�݊�=1^��U�z�#�ͱζ��:���^lKcw<�4B�f�E��hA�*�Ѵq\w1h�kuL&�,�s�~~<�b�%�I: �훖��r4]�u�PX~`p�����dO81�1��c�K�M�V.��,q�,�q�N��������wQ��K����
��ۚ��fb�(�Kb��$�j4(����d�J5� ������Î���㿟6���%�lQF�%�Ȳ��CїݚK�A��P���@>�����Z��w��I5��ӎ7Eg�v�|�N���Y�H\	C�x�E=�#��zD
o�@�����h�qx�Z/j�d\���~����
��,��ԶT gzޝ��_�`_G<k�O�R:�W���H��Ќ�n��I���;�$]��$P�BN.iU Ֆd��}�ᷪ���t�y�J>�ވ�uD�4�.w�B����<qm4��4���*f���X�пf������lf�����Od&�%p�|��:�8&��!ke� Ғ���d�k>�#r�#ֳ֚χz��bt2v�K�Y:N����Sī�����V4��Em=����uQI>m�����k��He*�>x�-�p�� 4F�Y�&k�)S婙����s`d�!$����~҂A�"[p���Q0@��o�KѸ^�Bئ��Cm;Cyt�+5����s¤0^谪9j­p�1�C��
�}ʙ�w��w���D��-\��+o��oQ�O1})�~�n�u�;Y��2X��$r�`���t��
�N*�������pQla˫x���O�R՘/C82\��Z��9�����aǴF�2�Y,U��V/� ��X�qRJ�L�k�R.�^��2UQ
����z�J�	�F���R���a>hd�/.�����0��4��p��U����-Kb�#���61PH��� mZ#V�H���%׊H&=/Q*H�b�Q��⦨.�el�a����B��n���Z��f�(~x�`�'�7y{���]v��#Ս���Na���5"�y�>��F�HR!#0�Q�/�w{A�t�Kdp+hZ���.&��?��>�1��>܈g�tr�q��(��f���WU�e�A0 �>	5���&������Z��׸��i���@���(_i���l� ��k�j���_~ �(��k���{��]tmh���v�@6��l��҃�>$xgo1�o�A?�|�܈��i�\�z:�yi'�)�_-���i�9���Ɂ�o�3H=V�3֙v���i��Z��j����/��"�+3g�KY]�If/���1�7�.V�ce��tx�D	eH���MM
�P230������e��u���ns��P�q�� ��d+���<�\V�4G��"���E�l�
Y��H�ֈ�{x�w|���4ۙE s9{���b��t���y%��Y.�%zk])��iuG'���r�0�و<�=���9	�G�cۘ��_�g�?��g-؍��H�9xt�.��0{�s*�G����'ޕ`�<�*'v���,�	y|P<۸N\��nFB+S��C�`9�>)������4�ظ�P2�;U�OX����t�� ����	�1�
ْ�t��`b�TFj#��u���f@�����j~a�1V�j�4/��Q����0n�;Z7��$ds�}�R����{�ƍL�� '>vf+O��[�يGjqZ��D[]�����4��(P d�Y�TMj�	�I�;"�@�������Xf��^C޲g�x0�7����x�A�Cd������S��崠g����0z�KC�[�pjz|���2�=_6���������jK��Yԇa_�}@1�f`2�9�Z�v��	�I�Y:���oXM������C.�_�NĮ�����L�*=��]�rkͩ��9�[�,VP���d���Vb��
�A��!,f%�2�,ϋW��t��c̗3mA���E�	-"�&�oՆ�g~N��nq.�c��4�� _5lnCd��x8��a��5"걢�B�'ph��}W�',�k�0��v0��RA��<lA̡O�F/�ŉ;6�����9�>9Z�$\%���p<��c��ێw-�^.OE��Og4.�}T�qL��eaa����T�0+�뱭N3�}�v�cW��@�thr��,�b�G�l�F� ����$1 !�I9H@x^`A4Z�M�^;�<�rg��bE����6Co'�~rVi�Q��l� zF?8Mw�>q	k��	�ZC!/t��>���~`��ަ�����!<
�Ere)��o�(�E��]���	@�5Q��~T�}��>�<4E�ny��k|%��n-ngs٤?s�"�:É�L�M؟���6*��Õ����q�9��q���ڼ��;߱s��$�O�YN�0���g�ӚK�^&V�"t�攣\�E�eK��q��bŲrK���&�}�_�_�S�\8P�����R���`Q9��rmpD��j�����1J���D�L��E.JH�È������B?=�^��<����0\"�d�w'��L����6r�G�A��b~U.i��j"RXmh�͓b!p��OC��U�����t��G��w�E�<�j	j��� �H@��\Q�nW����#o��� gǸ���gR��xX�3�k�M���_�j���`Y��O�VjA�&��o��n-(MA
��[�cd��&u�����<�/�P���p���� ?N4#�dvW��S[SKCߊ��n�$�K�:3FwWH�@(�g���ߗa��Igw3��p���vL�z��Ea~6�e'�N��<ΨJ�e�8*heu�jT����}A�/�,L���������Y4���Q���� �݀'�{
�:����Q��S,�1��)�[�.Ӌ1�O)��(���G�	�$Ӟ�Et�����$�vZ�e���?2�i:sh?����/���E�q08�� k��l-N�4k�6����M�t�h��8��D���v%^0U�]��(͉��
{b���c���wL�����r��~`;Wj���)�1��t0��X( ���D�\g�Hr7A�zn=���=F��l.��IGY��������Y��ДY�@6�Q0-��Ķ!`�jm�]d�-�(�:�:6e��� 0�O�i�{�+X�o�����ڵ�H��<z]&��-mlrބC�.1^t(h.�bĚi�p�p �q�'I�,�G|�I��)3jP�d�D��vÀ����]��:��j^W�nl��	��(�(��qNX6��>φbXx2��i:cR{z����>�_�+ϏO����9��d}=�cL_�=���y�$���߻UUB��W]�JC/`J���#�G�IZ<{����a���u��\9�>%�F������睚�g�(�� �1����<
�iF���%+\?3u�񱃊���tּ����^��X�����B����
��!���Uz>�1;�l@/W��d�b(w�n�2�4�H� f�&��-����Q��r��܏p�*�$�e�#��\��2]h���8�P���"�q�\M��P ��;F���'|Q�4ouvl(y8��f�UB�	�|_��'��o� #�)��&�@$�����^��x3�qNU/ A5O���ķ�(3P��UBei�ou5b���Y��_#4�(��rv������&o��7���T�3����e����u}�p�0^�&E�����u����H�L�����$.u���H3��k�+.&V�%����5����58���?�3�-���9������)T,M�9_H�`����N�V˥�y.T���T&?ҡ��{2�5a��*,D-I&���=�:��|)�9��j���dt�2V��Eq0�w�6�(�%�@^�ܳ�������;��O�ܦrmH��	��l=��Ox֢u}Ulg�������=ٌ���=�d�0�O�LV��[��$y�n7 s�ﵚ���0�;��\5�G+��(��t�����1Q_���aG��kQ��#�����@��R��BTb��J㪧-��?i����1���͌���τ(aܮ�m �E�lȤ
_�R������2�_	����\��Ks��b�Cr�y������c4\�`�Sj�A8�h�	E��&�5' ��чg���$�puئ���G��V[��c�D	�ZY��x�Ù���Һ�+�2ax�j�	��(��A���dW:�ƹ?#���B(�ؙ�oˬ���k	�bޥc�/*|���h��\��ʁ,5�*��Q�U�C�5�޳�g8>�^-��-�֣�1�ۆ0���1����Z �C����u�����ǟ�6�9��0UK�k��&G��S����p������n�!��Páh�DQStP9A��^-e�{t�H�5+>�j��l�����B���]po�*�g���%����EO�W�%-G�1�5��)^�(�0��f탠�v]������_�O�hAe2�GĄ��0o��S�	��6%祙�i��<٣��`ţ���QW���V�E�����[��96�6G�)��E/Qe�y��\oQ�[�#���f�Ffl^AX����~0p�������g�K�cQdgF\��q�x$P���"��� =ej	:�Z�r��m���"[�U�W�{6�wU�d^7�.]hi3ޝƀHbH���yТN�!#���[�j�0ϸ�C�@��AZ�����ڇW5�yq���$��Ev��o���n������-껳_���]:X�.��m���,�8��"O�����P=<^Vi��A�r��Qxv�y2?�L���B�O���	�Y�"M.� �Y�]�rSmE������ZjD����62&m#E�[+ J]y��-�@w�sfG��oov2���QgPƳS��8Gˬ�ko_ݩ���--P��GS����P���1�� ,�վ��Bc�+�@s�i�����_E�G�'b�����$���Al����2��`~���7á�+Qʥ5�F������b����C;)��|�p ��w�	x�$���Դ�a�R2���wk$3w͇1�^Q�&�,O9��^�>��.��[g�H�W��F�iYc�eWM�7dN�.������6��7�EX����N�L$�.g�Q� æ��
�����;���:ٻY�s���9#����*�&92UZ�Z��S��9�R{_��P&��	�O/v<�N���3R���G9�ͳ���Ծ��]�����&�`��u?��ᒈQwe�yo�����L5􁺪�U�D̅/�� ��yɔ��R�[ "��z��:�b32��1�Ѓ�I<<v/)y��t>z�+���#bl����\emq�*˙r${�g�{�i���Y������oi*(�!QT�F�^� �В_f���B[�g������0�T�뒔��G./.��0�$���\K���׳n�=[�Zڤ(#�<�]�7�SH��8i��'�K�j����1������$��iy�����^��f�??HTz8�΋>��O��a^_��OS�Is�-��)L��E�������
��o�VJ�H���-�r�9����������W4/���Ŕ7���V\�%5�˃�2����5>�^�=Qm��G�� �n�O\Z�&���#m'�/[�Q�жx8+N �2v{�o:h�䡞��G^y����'�3�0(�h� rTL�	mhT빩2�^�Pv)���i��i�����.�3�w�:e2K�b��m5��W�&�-�N���ED����hwo d6�U�tu�'4ݠ�`E噟^��X'�S�t����=���ƹ��������e�P�5�w��B	Owg/B�z̠�.@�8ȷ��!Wjk�G�w��d-���cn�✗���M�����{�4|`��A�=�ڥ����ב{j�v$�����z>�i�kwT���	|�o+F�k�Q�z�42�Zk1�M��e�㒾5��<6`w���Y�i)BVLh��Ǵ������V].�.,�x�����t��be��_�Y!oE���ح�Q�?�M�Q������K��xM���"F��:3`0����Ie�5�N���%��7&�v7����(��Q
���Z".U�ћ�&����O�""?)k`�?�C��o��(�s6H?�_�x{�q��8c�Ka�t}!yD�����v�j���e��_`������|��Wm����ѵ�[[�8q �/��F�1�%-�x���\�m���0�Jg ������)Ӟ��6v�pn������ϻfN�@��7��D;o�gw�<;�t:
a�������� (��{h��D;@j[(`�I��^ȱUf�75ǟ��lKѺ��-�Jd�
��m�%�
A��@�	.��t�WXM�&�9���|Cƒ(���V�TE>�  Y�kQ 0������"��E23%j�=�v���%KEe��� ��7�H��K��[*�jY~��8��8�*@��:�H�B;���U�ֲ���~FLR�0<�?|�F/������y��\�&c3���T��u˰�%�ҷ8a�l�ơ�`�$&z�f<=��&ZjCΝ�K[{��w�T�?Ux��G�gĖ@�v�?\9�+��vgq9��ި33y���
<���z�6���q,�[[X�Z��W}}"H	�K~+���۴?oV�$�	��΁<y�/-3�ѳ1"�Q�G��m+�<�dg�[�s*Y�}�\�iy��v��f`�����C}l�Y�i���U1��w5��I�(����fEGa��Jv'����	[��Z.��ϳ�ǳ�W�ڔ�Z{��ݝJ�|�t+���np�}8�4�C��N�?�mٜ�?@ʳ�I�CtU�R<��W�Vz=v0gl}��Zf��uq���x��-�$������6�jx;UPO�!�-������w�K�,���v�����e��)�
=�$�4r��0,X�o-!�f*�X7{r×�Nq1(�..��,�Y�t�GA̭���wǢ�$���3����m�=nĔ��O�RSD�2��	��:�����A��Ƭwav�vC;�c�,��X��2���,���l�.9:��B��D�X�Op��%1 �?}�Ɂ�߈b<Pe����Y:��Cn�.��G��o)Cͪ}�f�Y������0$P�g	o��x��wR���@D�A5�~�+�=�Z��<�r�� ��]��e9���fZ�6�id?���ʙX�,��D[ܾ��8����]X��H�?�;; Y�J��z̶��yD�<*���u�]�a�<Bc���l�	��(�-�~^��"��HQ{�H+�"*	v�U�Vt8�dxDz��Am|�9�]�5��G�(�Vd^Zǀh��4yo����Ԁ,Ny��h�f��0������ɧ�!k��;c���4IaOd�.{5Ǯ�* �&�K�B��h���q�A!���{t_�M*�hg��r9�%LOvmx�n���G	�$s���	E6���KrFg�g[�ha�aE�5��&)q@JE����<w�����:+]e���^Y�v�9�B���lh	M��.����q�;� ��5�����wiK�Rh��kj��QՕ�̽}��v�����Ƹ�_p��M�_��tWMr�p�UWN*r�ד:/G��$Uˏ%���e)k�뀉�e�q(|�QW��i�q���R�A3L�O
'��f�/��X�+���w��+��|4쯹"�(4W#�Zx,(S6�+���S���>G�96�#4c	 ]�$���,X�M��q6�t|���U�Mi�K�	}��?��B4b�>4oh�QB��H���O�.S���c�Rt�F��h�����ҀcM_�Sҿ|r����
mp�RX���ߜ�{@���0� �J����q�s4;�`#�H��n�ɾjn!ȵ�z�O��
D�P*A�{n�\܍�غ�D[Zu go=�"�~�\Dnռ�[3���E1�Ӱt[����Y.��Z�"�X�&ǚD�p���Q ��5��=��¥���[�iQvC��C$�vס>?ٲq��_�f�?-B`�R�[B�~V�htY�_�O��V.�	�	�Պ9�#�F��`���ņ���w�D���>47�E�b�����ݭ)��Y�^�4��s���	)*Ħeֹ����n�c�������:?R��&a��9����t>5^k �պ��3���!�2Q���K�MI�c%#�H�P�OIVh�>˄�N{���E�"�_�zL/P=5���yn*\����y=B��AHo�$č��%�Wl+BF������֙����:(��n�+��QIޠ�����2��!KW¡[2ֱ@��^N���|�|��-w��ݲ���v��\z6�,@a�=K� ��Y��#�{����@����lM�H�*�<�wR�'��e��(��zY�^�̵P�E���%
�f�{)-��* �0=�v����Qк��W�N���T~WXEz�Q�ݧ��
�%��R_ե�S���m2��L���`���0a� ����6C�r�C͗��|�D���mW�뿺��fu)��N̐����4-5`v`;
5��]G\��e'�s\�#vΡ����Ƽw��Rl���{��Ѧoqp�hB�́K:o�g7��guq�B�u�㹘��q���qppd@� ���ƙ�V9�/�0��ߴ��uv����180�k-��Aɟ.����Fªi٤�[d���e���>�_rcmT������[7b�kTl���qѹ�5=���Y�W-�Q,�1X�����1^>Â�i�	�o�����GeK|�@n��X��$�9�ԣ##�|\��	��t��� -k���=����
��e��m>�8���i�k�k� º���@�T GŘ;X!i�=�  ��;���vEÁ8reoq2OG�Iw�z��,�3��'$]��q67n� ID�@���]��z�w��4�%{����8�.vߦb��j�h�^\)8q�}���ԉ/����:���;�?J�g��b*�'���fp�{0*���RFؖ�hƤ�./��[�;�R�V�0b
-é3K��0�6�T!	����_��w�X�yjX����i���mO�7��)`[�%�ƍh-�X�C~��e�
;�g�CxD|`#N�� ��C1�X�|�^�7i�NwE*��N�]�TG�Y��}#�uE���f��O�:�Fd�Gvm����_R�{�A�Y��z���X�D��T�E�༃��StsCS�"�
�_���J�r�Iհ�S��!֦�!������ƀ7H� ՟sҙa}d��Į�l+�f-�%?���`8� �;Wn5B�DR��G�r�1��/h�2�"�͜�"n��h��z�����sH/�5ۆ��g!i�E��(��6YC�;>Y���pz6�_w�#�W���s�c�d4�,�}u��0�����7R��G?WҼg��}�,xgp
�ϼn�P�ķ~��p{o;��Ӕx�x���x�
���vʴ#�9��k�ɥ�Zv>=��U��ˢ)<��� 9ΐ�I�ӹ)��<.��`2����a2W6�KA�W�}�f-ϝ���q��p�O��r���+�N�*6Fh��Y�+r](𤨷�A�K�b��ٳ��t���{��M�h�m�6z�#���_QF
2�?^��+��jg�������3��1T6;(�!��$b=3~�H[[�pf�nJ=�G�#,dP4����Q�E���y�^P�����9�.�ғ�?rMꕢJ$j+E����2�Q�?i��:���fv��|r�AZy�q�~��i��,�������]���X�u���%0YZr����?���8[�r>� ��;�96V+��ܸ��h�k�:Ӆ>j���;tp4sр����5��q��d�m�m_(5����`A��Sn)o$��U�4̲�KG=ӛc�������K�W1;��%�52bp/�"��ʭTq�3�A�z�^��&WN�w�Y�*4߀�M�A�8VM��/^�%P��pɈ��K��	T��	�?�5v�~GQ����>�FQ���C�/�l�!y:l���}���j��qQ���J��8�G�[���oQ��MZ���3lF��؁S�0Qp��-l��d����8Ё��/�q���Q��T�di��t�������ʼyH��|���5�/��\4ϫ�/�]܉���-�np����������� -Ң����*�k�#5K3'/i�@�ͨ�F��g��[S��N�<�s5&�e�pa�����j�?�7�4�0=1c0�L�C�m�в'�W���m�7��tz�T�:���r|���IǊP�z:������^ �@.ɮ!��;�
���a�^��[�n0p����3����3�ɷ�xX�We�J����f���{��x��k'�T�܉�zx1i;�D oR}�����������F�o]a����6�=^���8s�0��ȣj�ࣛ���O�\�v5T)���7�rL�U����+0;��g���:^-0��F��
H�~|�jw#h8�1��!��/W�>�k�6�o��č|Ѻ�HQ���6�˄�)���dZ�@�d�GN��aT/�t��F���8�T�ꚳ�\AI����]/�S��V�r?	~W*���h2�u~�7A�,�UO.ٜ�a���w��}�@D�gmˌq�+�;�.m�����)[��V@�S�M�f|J1��u��e3dղr�&A��3O�f+�}=]"��RGJ��G�/Qڹ����v�P�[S�;�S���݀�󰭸s*~�Z�$��?�wo�Qz�h�X%,i�����wf�ޔ.�-c������	���T�9��v��J@���Ҵō����SX�����]��� ���<������Ax���Ӯf	 �ap|���>�dX�����FyG��?���-<QP�F��f��hO@�!�����sd9a������ �6d�h��hT�[��܅�ݷ�Zu;	���G��c�E�y���C���ZQH���R��2�29g81��!9d�ϥ5�|EH�B��/��R�!��i����IV�su��ڇ�����u b�
`�"5�.�*�֎�%G�_���ߖ�E"G�$hc�1O�2�Iؽ��1�����C�S�
��@��?�"Oo�t'�e��(��t��*v�<	�Z��!�?�%b�p���
�/=3��)��I#%tH,��J<�M����>�'�W�/8���]��?�riE:gi�< ��
2���M���^[�IF�ֹ�T��\�	a1=K�P���O�3�l`�I���*��@��+�8���s;I+�>}��Чv(�@���|�}��~��(�Ld�]%�в6�g��*`Q������p�k� �.�N�|��$pr'b?��K��p�lg`Ji���w;P\� ���j�&��i�Jr��`_X1�fӼbN;�����v��:�B�u�@�y�T�ο����e�ly3z���+84�V�U5黰�{ă �>ìws�I�r�I���.{�6��Ȝd2��UD!��Ve�����ZĪ� W!_8���Fo��)7Nq>}E+�1����A���9��v�%��@�&Fp��0�(������ne}B��P���.��g��˴u��k�pR
���Ddb�|��Fd��W���F�\hlt��f�
Oxj��F��dd��J�[���Έ�`=�)���ݲQ/�� K�f�]Lũ�.RT�Y��u9w�8)9�k%\ꐢrA�0��8HЉ�d�؆��\u��f�*�ED]�}]�g -�I�=ʹ�ܻ�x�u��.`s�!5DyQ,6�]�+�"����Ƿ}%���<���
�:V�	��ǂ�@R�>o��4k"@�y2,��˲�ϭ�uB18�q=-��&�d쩏�?�6}� ��IS�2�:bGV��¶L�:^ �a��^U���^wفS���S����� �J�$\{��!b]4D�z��Vu����<R�u�5����-����8t[gP�����H��YZ����0�z�mP�����M��Mx��+��?#a�h��A�X��h�_4�% g6u��y&���
��s��L�
���i��-^������yZMY�=�&����{'|,������ԑ��M�{˯53�d�k�� D7]�2^�2:���u�V>Z�?42�(^��11��<S��ۧ�v"��Q{%w���3F�����RG�E I�%�����jq��~���۬פ<��S$�*r���&�M���ۜԇ��4��ZPg�$C��r9����������|_�Hwnk�? ȵ���r��/����p��f���k�WH��
����|f�D�;�;��~�L��I��okl�^\l�(�� ��s� �4���{P�,�VX�i糶�^"���v
�G̿,�q��t
��~��˱VB���2�Qg���s�}~�0P������J�"X*[�Nث/*�����D�ϻo�S��zEp.m�B�R*@�.'j�}%�q�u�I�2m��+�m�!f�={R9o�s��|[?���,Y�Ặ���c��.����n-%��V�i!���V�~��[@Pˊ�*(e�ǯ�ƍ۲��A��WT������{o���:'/�)����%�݌.v���#P� 	;80S�8��ͫ�J�ݩ���M��1k
Y���j{�^�~yq>?zg�Y��)+��my�0����jnl�`�[<����W7u�<����<��6֤��x�m�e����<��-�� �^1ҡ>D��3�U@��c�h3�.�P�+z$/B�ᱢ���<Qś[j�	!��W�2�Oϼ��=�x�:%�Р�3Lr3�_�h�D}}Wh=S
��:&<�Mu٩�/1�j}��~��Щ%V�,��vE����bs�7^,��]ꓟ�nڦ�Pv��B�~X��'��J	���%�X�� �FH���Q�����ds" ����C7������DZ9�"	Te��W D&�Y��}�Aޓ�w��;��/H��5l��[)]�gQ�82s�ٜe���\�eP�|���C�˔�А��2 $���u;���hޘ���xվI�O���ٯ��f$�$Emiƹ�QJG�{���`�,�b����.vL�H�}L��p��~��}n�Y��pF'a�S	4�'����;	B�x�	Rz���|Hy����r��ʜ�@����l�����(�g�J���J���/9[��r�џ��U�
�a��wC�X��q`�-�� �@A��-뗯Yb�L��~ї˹�M�X����en�e
4T	��`�����8��KZ���튥�����3��P0���c�P���3�A�9L��cL�u�a��~D�\�_��g;���銉�<X������OS��$�HC#ʽ� B�/o���1��&m�W��`�Ĝ���8�𷟵��R1��~Ɗj���������L���\~�U�0`���/{H�o7D<�H뢵Cv4Ki�҅-^$����ϋ�]�γ*�t�O�����?��K���9�w���׫��NɛT��&h�DW����y b�GB��L��)���\�����g��^�R$ED"t�,����+�ʓ|��7T�W�B�;(�#���"��Dֈt��S �I��r��\Ŝ�����w��;��J��3�BAt���T/��]dG�2�| 7KH�9�Y��|.Y�C�������n/��o���t����EZ�3�^Ӝ��x�j��npD`�B�"5��,�-�Rbހ�.-Y��ݱ����uO�x%��qd����K^�z��������N��xo<��c�N��ػ�ܝ��w_y\蒣��s�"�캇���i0Ȉ�-t�9�d{y���������!�_�;�tT�}~�}.�͑��+�Խ�<�����v���y���C =B?����Z'�a��{�/���@�4�K,9�t˝!edA���B.W+8��٠�%7;k��|z	p�1=#v�2˺��1�f������
8c�}�V��������'����xY��Lw��I/�$�P��B���]�3S�^U�Xȡ��	��.��Էѐ`���4����2����)3��<�=�<���ڕ�}�?�=�
��Y����BJi���a17Q���~G}�{K�P�%u|�O�M�=꧂�6��K�yVXM	�]̞) )�e�͂.���)�dMa$�!���9i�	85�������i0i{QL{�:���Q���?&�k��> C,�wӏ�d��?�s!���k�z�`�}�n�������YFV*Lս3�9�V-qE��dB*E�}�i�6��DJu]��1���+ N�+>%��/wj�	$Du��u�}�_�T���iN��yQ���[hQ+7�C��Ж�̄K���6F%_9}5�(��Q�=�j��j���RX}����ܺHa�h��f_����s�]9*@�����'��p�rg��\�<�������uw9g�y��K��C䇒��~�'�x�'��+1r����e�6l]�f�`�9i��� 'c�3��۷���h��x/~&��`�Gd$�T%�ס�$<GA���O]s�ry�齆#�-��;1s���@s�秥����
��m ��Дlʟ����l�-d��tw.��#��eNm,�dU
��5���v}�_�H���n"#X�b��n5����|yޠ���*ea�Íjv�'2ճ�nt�h�r4.��|��c^�8�� ���o	�2N��/��e�7ёi���\�l�v�[�/�,��s�k�s|�$�AW��d��
p"���ZA���1�?`}v<C��:�|����4�;���m��~�e����o��fċ$�CP�g*o�A�d�)i�_z@t�H{��i��F"ת�!6��r3_��H��[��:3��Ljo�v���6X�Z�ZZm�?擀7�ZA2����ĸ�|�M�l�?N�F=�n�J�w�r�{"��1��sS�y�׳�]T��T��~�V!Qhk���۴�e厀S������w����ƈ㥨=�d~�0x�ɛVnZ�2������a��u��f�������o~W�ͻ8e�
lx'+:��[���Tq&)���sD&+u�﯊+��˔!��qO�^�Z�n��lL�u^_����m����a��X�����Mw��D�lƇ��N��2v��iv�YVk�2�Ni���kyiR����2[I5� �AX�<jA�RZ{�w�	ٔ�NT��'�e�T�IlM2�#E�܋�V�+6�"MFd[������ҍ9}�v�����#y�����Mzy����<k�c¼ug�J�a��
���,T�
��)��Q��"e�qnirS�ֆМ�Գ!&
�ܕ�N��Ǖ"5'�A��q��k�F[�
�<μ(+8'���_/�b�jF����%�l3�Rq<�>	��P邚����v\h��TL��7[�S=#��`!Ѣ_a��8�Y��yR��HK�t:����~��3GU�����j؞����.���?5��]}`b���?3��6g�?����������+��X�쒘CU�l��}p��~6�gR�SØ~ 涜��������_1}�.���mHWd&�_ʺ7�N�w�T��y֒k�<A�ɺW&.g�`��k�9�}" W�� )N���PwdA�S$#~��i�+�G��;�OZnk5�W:�(f�;"�B�Il��{�vE���"�'�rb��P�Ux4Ia+t*H1�y�%��kO���59Q�#�V����?�'R�?�o�C�w�Y*5��$��:y�Z���:3bi1<Xb-}��r�ޥ�����wC����^Z������4(\R�Bؙ�͍�t�>s�"���v��O��]����'�����(��!$� ����~k�Y��I���Q�W'nţU�mq��Aq�V�nmE�G���~��Imaj���P�d��M��W�_j;���H ��[A�k@i|��y\Ư~�=q2��xC'��u��s϶=�`@�~2�Qy�U}�p���"���㧇��G�=��EF ұ�
���@��a���4�uo��g�[f��o���b������Κi������D��� cɨȊ̓'�hH%5�{�ʜ��rt�{Ml4��L#W�K�������	�p����̟�,����, G��בL\, y_j^��n=���1ۇN��"zpkn*S��D;
G�gg�����
J��m7�`ɉ��ސ|�G��P���\3 �f�+�9U��JI!�" �U��^.������b��6�&��rL�P~��� X��
T ���C�˄z��w�v`@n����ߩa�6҇���g���obRU!���(_c��9�{��b$7�܉���F��ﰴ	����uh~�����pR��sr-����p3�����՛��y��P����ѻ��ά�d`bW)���j_�Y��{k���{��yH]Ӱ�xކo���ac�s�X�N}	d�[{�a)������\ڞ$D�-�W�x��N��,Y��\�f�ߣ�ڑ���J��u0�?RW���Ѽ4�Ax�煂}�s�3wER2�:��Ǚ����T���f�-�<P�Z����&�ag柱AT��t:��~�2��x8�@I�RZ�7}{�,=��V�0hؒ�y�6�=&/b�k��#�.�D�?���`Ck���W���q2?��KY�%�2��xs���o��.�b��܃�)�xn�=�RinU_�Ks�����0��;x#7��)C�76��UK����*wh&���x1����β�C>����A��WuSe��k�_&�܈;�[�:x����WJ�Jf��4]��\qJ��U��aO����5�	�X}��攸zڃJ�\SW�}�����`�xl�%LxZ���Ăv2B�:�r�1.�k�#�M.������I(�D�I�Y*�����:�>���F���s���K���7e9�$����ꤳ&ֿf� ;àču��J���o�<4ѓ��� q��fX/�Ɉ��F�M�Zl���yo
��a�g
Y��I�CS� Q��b�� �ɽ6=�J�ƛ+��!��0�5WL��uj���or�Ʊ��[��[��gްjE^틈Dx��!�XC� cl�Ҍu�ԧi�#څ���^���O���x�	G��_ܩ0^�6���4}S��-n�C4'�`�Ǫ}1(�����q���?�	c�)�_�<��d�j�@ҙ?~�)��j�RE���b�[��h�ɹV�>�b~�
�z�m�������QL�Ņ��K-8���Fme|�$�RLHĈ�L�],�����Od{�'��X���P�@�9K��ؕf�fS�^���H�2���6�#�a���B?W
���9$���7|����0-�h\��[I2Np����=
���A��9u|m��"B�M[�*�C̗!�/7���SV&�;͛�[�]1oA����4uW����F>/��W�{ �n��/�p���O�^pb���2cq5n�+�Z$[�J8��O!����	h��޳���8�9K�\zf&,1�4��r�\f�-�ḙJJ+m8�Iĝ�8�<�0@K����� ���+�T�!��5b¼	����\;K@�X�ps1jB�I�;���<
�H^����w��<��a����1M15��p�l�CzƤ �d|�A��"�6��I���:�H�{+ȋ�8+nb�qw'�Zt���_��|ge�}i���H��������Q��,����q��G�����+���<8l7���<=���Pn���`�0#:��Z �&� 9mc�߇�L��z��<����"X�
?P6C6�/=q ɝ���Qx��㪌��#�P�֬�{˷�Ov�ş�I�K@F��ǯ�=�Fj�"��.�Mto-M�y�Z%��h$ ���Y�Ǥ|��f1Q�8�z�&�� �?�5
�'�a�\��gc���J�@o������`����rT#(6q��jcM�\�
OR�愚O^�Ѝ�/���Ә��m�A�ϨXK�*�y�%�2*�Q�J �sK������"F�B�V�$(Z��ӳZ��¦��j����UTi�m�!��� &�Ȗ��Gp��;�_�	�)8��lK�F���z���}�-��sw������[/�[��@�(�ի�'����a��8�8v?��{ �5�#�� �Y�b��y��JnK�z���}{S�J�s�f���}���� ,}�-vq����Kk������L&�;wM�)�t��t�J/�$������'����T������%��ϸ9�th 'l�D�8�e	R��s(���Qt3���["&�e�MGr���&���w�d�h_9�H��MS���Rd}��X
�U��2�r���rq��Ga~�H��#.RW��M����N7��a�&d�����G��3��T��9Y|d.0A�@�|Z�Ԡh*\Q��1�l`�e�L�
���b���p�)�)���<��d����("J�t����e�ʙ4K�� ����s���0�R~��e�UFw�:��O9u͹E�W�SFL���u9iΧ�2cRc��w\k�[�@�MV�d<l����|�8�R=Ȉ�L�`�/c���R�u�z�ݎ�{(�1&��+�����\�~i�F������d��]���)���(����騰��m6�Ķ��'p�7�vy&��	���2Ql8�j�N�\�C�g�C�����/M�peLn�7�:����G��7m�c��E�jAd���Am�10Z�S{@�� ��˧�ƿ�p�JUZn�_���.>e����l9g裋�,9DE�0ڀ`꣊���+	o!�޹+����LZ���PO�%µ_����K �T���e��}� ����^mG�O ~����s��R�5�`2�>4ylk�9��9o���膕�ʇ����L���+���p�M�̡�U��B�M��B��M�+؞�۲���ݨ���>Xg!�f�/[]'~ՄZhV>�[��9��5�W���@�k��ե\�*S�(���h���-*@>8f}4>��vjo�9Ӱ��eV�	C��t�"%@��2Z�,��b��l��Ћ���Z��$`���������y���<����Akz�{!&�'41b��&o�-��w���C&�b�-��]��U/"����gZ 8a��I�J�-%L �hւD��x�ȓ�ׯ+�<)������Su
�>2r�!~L�4mi*�:g�b�M���ລL�c B6"���7���.�;�m0	^���
����(|P���{��]�;�ίߣ�䍹��aU���r]�������R�W#;?G@3Ԁ�-�Y�|�n8����8��G�,��a�̣Y�WƠ�=PTK��\UM��t�,^��h��4�Zr�H��t�+s��:P��j�gU�@A�M����G8;
��I`lԬ�?�%�M�l-n0J$k*#4R�&��m�W܉�ϔ��h��T9��Sk{/&�X�`a�b��t�}0i��^r�z��/�/�1K��c867��1�A�-�Ai!_8�hB����7e����=�\�-%�PzN��	#�KL�[���;�C{�E�0!@�~�!r���D>z.�?�̚>��Iq������j����:k�R��x4�D����LX�����q,ր��~#�}�MV���
�#�����¿;�Nv���:��e�8�*e�+���>��QJ��ڱ�ԬS��l��[@l��]��ru�3��w$��M������2m�b6j3�p���6ԯ�$��%���/��z,�fXR,.0����Kr��q8-���o��>��I�fe�E:_�l�NpZ�8�,+�SS��ڎ��;T�n�C[���)�
*�\�R���������
ڸ��ܑ0Ұ�6�t��.S|����N�HR���W��}�_�u*�U�_l�2��ℹU4v�y��V�,X�V75���҈^)}��Jb�^�!��͢k��g��S�� {�,؀�bA���}x�[�����1'l]0"*���jv�� �"���<.��5��'Vʶ<��ߎ�@���D�;�V��LǄt�@F� bk�|�c�ō��v��Â^Y���w>�^0��.�����^a��.����j�r��%��a�V\pi~��1�	����Ź��r'ۑ<�z����_�6û^�����#v� ��Kt������7#R�-��pD}�?�0[��ܢ>�NX�!F�*�9G���\Bjf��^�"����1��Ƽq[��$�S���oHx��ry5m�eZ�5�_"�9&�<T�e&�SoA��E�o�ksђ7ЄjL6���P]�K�Y~*r	�,�ȂC�ݖYe����<duM���%hr�^H �p��OW���5.�FH���WO#�۟QBE?����_��Nۭ�|b��ؚ_J�_���A�xx�8j6���<��`��}�D��i��"�GVxZ}������� ��1²'��j�ݘ��<aQ�Fo-���>\��Z�+�B�#� ���th�0�bV�3��~E+� s/o{d��S�"�/��}�,�7�5D�J-1-��	����NKD^ʿ�_/1IV?:�����rj�Upn �T4�Nn�翑G� �{��ՉL��$N^{uG"�(�`��J��
ۃ-���
�ʤ�7��%��M�V�G9�3UGc��NU��iF��q7Ţ)��������[����F��޶�+QtOꩯ�PB�$%g��#g��#"������$J�48��{�������{���-0��%Q 9r�XO�y��ۑ����!9wY\����K���� JEu��4ףGऩX�j�ⱼX�,�[S�0f@8��~1�9�D?_�VL:^�L}]03~��7:�c}�m	h������WJ}���h� U�%/w��	?:JF�.f������7$v���j�c���PX��22AKu�?�P�$b�A��}�V�F��E��MK�D2���A�=��n���Xc�)2%�py�������l[�wJu0T�B��z�"}r�g��!��M��=�ZL���Oǖ�if�gý)Bp0:YxD0ph�v�
Ha�؎ܨ@EK9 �i���R�������ǂ��������C��@|I�j��A�z�e�%8�x����wI�k�@�'�M��9���+��f�?/����{��@.��9�d�0j�f�@A@e�n�ėpI�p���+LzD��&��j5p{W-O��rя1N|��iʸ��Q)a��z��,W�=s1�͜�]�� 	:;��(q;��~l�ѓ�	9���~;9l�R�.1�X���Gy��ۖ����ܑ-���o-�%�m�N�l� �l5Q���$B�Y�"e���,�t�t� c[1���J�X]@U9J��(�kx:���~5����n�OB��E��s�.�T�L�?�\Q�iTV�p�/'#������~�y���q����u��CTf�k�لM؉��@G0A�C]6�X}�%�B7�~B��i+J��+?����ǇX<.���6p��K��6�0o��+�ЗsN�,'�l�8��K����ͼ֋𣫋+x��Jԑ��;P���z���ŝZk��aI�I��6	a0��2�I�H��,|�\r����X��f�5��ץ�T�Ѡ0���GƎ�2�A*��|r֢�B�"r�f"A�G�b�R��O�g���w�ò�,X.�/�:����4�����$ri'��Vn�?������f��+���Z^�n�X��k���p�����_����bG19��E� �G��Ӎ�0n��S���,�a�Ե+�J���mZ�ʱ�ǚX�yV̆��"` ������@pT�+�b��/!������|�$�]��o�0s�ɓu���ջ��i��������0ErU٠�d?���s�[3(���َp��G�z�xc٘i����e{iF���)��,a�}�>�ITK����;�U��F0؂йXNQtVC��0B_��p�̎\f�,�WK�V1�R?⌒���X��|��w~�&�� y٘O����k��pvy獏h&Ò_;�N��s��K�?�$⡊�e�D���@Y1�t�5G�򑟘,r��U�?��5�>�GB矟��`�r���!�+�%:v)��N.�b��	`5ީ�g���f�=��QMIz�V��A�R:�������6&У���{�,sy� �sW���C��`�@l�>A�O3^�KI#���cY7��� ��lnx2�"ⵎ��[p�G�����)��2����`U/�a���,>�{i[���+�ǽ�p�D����H��D k��6T!��
����6��o�Ë?"Y��y��Pw1��HDE�TyI�`��<o���d�OVyD�98�5W����,��4G��cq�|D��+�tf�S ��$ͯ *!�|Js�z�� G�u&l�����f�,͋�7�bxhx6~i�g�U5N�G��K�m̛X<�o4�j��~��b�ZΤ��(��;�2^���u9���p��3r���x�~��§������{�|Fv,��q]����I|�zXX�l�L��>P�(,�(��ts)- �4�t�g^#aȃ%r �z������Sm�i]s�@�B&fr��O�R	F�U�gj�I�y�$�}�z�����?\*��G�׵�#�]�1[�cM�N�T�O.��2��V2�&�~B&���q`az��r9Z��x���|+��f��o�OP�62�U�Y�Jv'�4�Sn����N�֓TL�fz
:�xDR���L�qwb�1�$3����`�j���@ӛ 2��ȼ�L�i��C#������QH�Q%� 4z/�t:_�y����ku�'��Uu��:���ㅑ�G4���v�[�Ό̳�&�!Q�9΃��d����u��^8	Y{��M$ǁ�Q4m	�����J�w����rT���!GN�-K��;�G�\#uGӻ��Pϻp#�ke�,ǅ?��C������1l��<4�:�����%J3�Q��������V;���uď?�kx�첗�z*+�D����E�_�W��bN:х�7��@nOY�y��~��Q��/|��Y�k�����tK�H�����Pj/a�͋b�M��r��(4U���Rn��LZ�x��J��w?�M�˙ �q'�|$8�0��X-:8�g("Zks�1�.eΗC_��2�A�
����l�X��.O�L�v��z��a��;�wƛ�
7�K��<�֩�`�{Y�<D�&�P��|��`�t�$�!qe�}y����
RA��{�4F�0P���oˢ��&TȐ��$�s�M��k�=T�bcM�k��09�Ϊ�uL�o�uA۸V�
+�y�=�IUʌ*��D�l��K�9�:i�7yx�	'K�5���~��W�PsQ���nRY��w��k��l�?���H���~�@M�����h&D�k�9��R־��qUz��.hwuG��Y�O�/���`"���h]դ�����ˉo�vjY��_�~q��F�Z�$��WM>���9u�F"��Tv��ݹ��De�tz���1��p����������Bb�`7]@iz�t�!�M�m+��w����q��h`2��9��:=ˡ�Pŏ��.����b�@H���,��X�Z�������4��	�NE��I��_,{�*
>ë�[�H��>pVD���tE	���"�ܬ흕r��B�ngf��D�I��O>��L�{;>���'ʍS�7���*>���8�V�E�
�#/z�>����0�2z�ǚ���b�@Z�)�cui�{v���*>p�hG }	͈"͔��G��[�2�mب�BW�kKN2�D�"��D�:;������禗qz��6���D����Zn8j �nlVQ�ܝ���&�; ���}��AܩY���+D;�������St;�g\{n]�B��#�|���i���͛8M�ko�Jƹ��s;����V�U��X���\��@�=�Jᯆ7�=H�3i��03RPcɔٗ�r���a"6���Ǜ�'���������b�����ʱf�e[��M�S&�K���Aە�	�,[{�ٱ��=6?ev�Kv[XZ_�}�
�T������ �x�]�R�����*m6���^<Ț��e�_�2��6�z^����hDf�1<=pj���y�aT���.�{�'NV(?�r�u0�#Q!��4#�5�$�mL��.G+��.����7E�kI�4�����sΝ��)Y�Fѵ�(�E�p�mN��֎ӵ^�m��" ��]2�^�=�^�g"�]�
����7���r+�)� 5�5�ʕ2x,Le
z����R��Rc���t6��wb��1�n��t?�.� v��~N��J1���;�?S�:��JR7�8���\|��?w*d��Û�qy3���΀L�Z>00�{����)*����Ĝ���"d}��xX�nٵ�����HM)�0�fK�[{�~�u��.N�@b����#FVI���~OTM��&r[Ē��_�Ǝ|x�I����:!,?�@���t	js������-���h��/ ��N�1a0�ka����&��f�!_�`l1��%�o�o|�GN
����_�u�t��]HKڽ���U�D��`�,�d�E������2(����~����k����k�7��� "�H��,l+��,-���T��6�0���x����]��f�D�!���ux
�)BxB`̋����w�S��Rw��ĉ͎|):|���Vf�˛�9>�&�ϣ��a��xЀ`:�����7������o��,pa2J{��|;���Vo�5��5mi�s���ꯏZ�s�o���Y�,��UǶY<'����w)r8�����U]ҋ��KlqA��\̗����E�ʮa�Srȫ ���?P("���o�]����I�*9�iA�O��q�k��}��~c;=�eg�p�2��z=)���ݡԦ�1���NA}k�L���i%+�Sͧ�`���!�o(�1w��>��@�v��`�ĉ��+�ZKZ���:�7�D�c�/Ս{<�`�x�k|)���łQMo��܂v*�ͫ���sx�f2BE�F-����,�.�[��J�Q�S�F[�p���'�J�ʯ�w�$yqd�V�� /�8W蔞�h��jW�mjQ�w`�)�gP|Q*�*�m�K�3��wהl��M��7ã|=�t��������)^	e7=��%��\����nt+"9�W�=��oX��bi���K4)g��� p�����zE_�OcдH�n�&:�yN�Y��R�p�U���fn�m}���Yu?�s;<b`�����jJS�L�����#t�yݮ�S�M�l�ʳ+�=XJ� +H�<��)4���oӪ�f&&�.7h�լoL�&����x8���r��[L�T>��t:��)[P�R)�1���Ӣ�oc�g ��	�����8��,[ӎi1'16`�cz�N�U.��}9�ߏ�	H�*�x�t��ϓ�i�U��/%֓^��(�q)iNus�x6h���ҏl}Z�h�pJ#©Vʬ��Q�>��78j���2��B�Ѿ��� - ���Ɔ��]��O��r�	V��HK_Pľ�����.06R��F�b6��k'���cO���_7Y�����}�J<���H����s��ֆU�� Z�#��:���ƾ5a�[�Аo�e���ZRܷ~t�2z�4n{����68��.Sb`?j�S���q��YBh�R��E-�� L;x�cB���c�@�SQ�p��\�2�g����%NgY$K�R%�!��/r�p�����⹂TG�G����������D��t�F�tNq�K����<�3�"8�z�Y�	5�P�nT�?�!�{e]�;h{V;�J
&���(���?����#�~ӱvÆe�����0��y�{�T�u���
��,���-���7h��̪�U��M4(�f�~qI�G�CL\s�i��Ҍ2�7=��p- �E�A�s�Z��IEO���gЅiD0��Q��}�a�,e�_e���'�� (_cqE�#W�O�>u����Sv�5���N�0�W@�����N�6��s�%쥐UU;'}]��$)]Xtl�|c����b.瘠N�;�`)-@:	�uG��,���R���t�7�G�/% ؓ���N5R����mq&\�_C�}4������ �O����}�LӲt�ho�%Dź��n�g�R�zjR-a"�2�}@���2�l��g�~{£��s�/CU��c�� �����0����<�����"9��1e,Y�@�L��$m���W��oQJ�@�֓@C�I����,���]ྣ��mC(�x�i��m� 
{Y:����O�4��kE��	c�
�[��w\�%�:ۓ�~�Tt4+�%�D�v��y�$��1��"��	�n@������«E��)�÷������_�	�M����L"�4��7��\�?Wָ�K��K��V���ї� ��_9<���lBEy�I��_��l6�zJ�y����]�
�m�!�!s�H�{�G�t,Z�g�iEI��^�
Y-��n)SS<\��=ذ[���Hs}.�h-��������z;��M�oS'gu�h�!����;Kd��I���+������i������D�|+�׳G��E'/����^�7�}����@�K�^�"gWrf	b�L}�N��\�p��m�P,�!�?Wjߎ�M�eP �媭)�\�]P�1"<u��:��i(�p���Y���B�١k}���.�:U�o�$����W��)�����}+�7���uJs\�nfiZ��Zwa(�D5[]s�k��Z�F}yn/"|ݍFC�" �;pWf'��S.N=o^�5���_��M�v���-	ݔ�{:�ۉcV�j	k���ҷ��������ٹu�R��a�x����xA3�h����6��?a�v:�؀S��5�1���u��1^�Z��nn���1��uu�2�Z�M���N�󭈔�f�QP}-�|`EĤ%%j���/xlQ?</�b*��&,-�aꓧe�~e��.>�|P�wWd����P���,rS���5CT5�i9�%E�\�p�)��i���~?��\��Q�r\]��� ��Q3G֌Q3^��d�ޜ�ѽ���G� ����!�r@��5@�����^{'�ibg'1���Nn��#)��=�ئ��f��Z�P��@"����ä�w�4�I��[T={�6D�-hX�z2*Vy3�"@:�_�e1&��h�a���s.������-ՉhW56��V�.E���(@Y���2kz�y�qPx�m�a�7�Y.�s(l;J�x�1�����Ҍ��,��}�	y)C�YHDj��P�`� i���=�#��o�7i�������I��]7~B���;Y�d�i�t���~}�zI����w�E����5���k&B���m��γ��Q$9�c�G,�I?��t�mWn<H���C&L*��_�zʏ!�$)[ ˨�3��]8��`{��z����y�ۙl� ������	̛\�'pM�)' �����N����Ԡ�o|b鰔7S; >ڽ`t�n���	Qz�|�eʛ��N�i��|��H�/}\�����.���n���Ȑ���a�q^�wO֢?�#�`��\l��L�l�-��r���د	bX�]�"����i��x�\9��o
�_��A�(�CJ�{�v,o:����X+$n��1(mnc/.�5��&Kw^C��V�Q����-�|�T��ߓ;����R���/"�4v��4=:c^��Т��g��DG3bXd�����w�{�%����>m?DI>}�+\�\J��OJ�$��P�6�V�C���c��~��<nד5�8�-K��݇���K�� -��.�������9����5���R������`�]���?�<8���"�A��v��3n�.�G���)/�(UO�a|hc�v�Sq�-�5�T%�ˠa�,mj�n�Ǯ��j�Ă�]�6���^ҥ������g)�}�
��4TW����V�ەh�w�x�BP�NM�AZxs�Zâ��t�]m��"�Pp���Gl�����/id����߂��>G �����G�ӈTS�d��q���uƾ������^qX�'�K�����X�ԘJ������=F�G-햰dz�|��[�`@U�\<KCkY��%2x~r�y}��<���Q1�ƿ�����I�郱C=�
�SS���r��#�5�yj˫�g�2C���T�1Pz�W�n���@��OMVjP;?���*L�N��kR��`���/�ƥ����0w*�I���>W�L�}�x�.s��j�d�t�P��"v翪F��>t���r�&�25�WN��{��o]�c���}R�1Y��3mZ::r�����o�~��Z"��l �1����������J�1�w��A��#��0ӛ;١&�����7d9�ڇ5d��b�`P�A�Is��U�i�UVy��^�W�N�1>��1�ِR�����A��A�`oT�`(�	���Hp!���D��\/�W��_��1�v,�ʭ�ʊ���I���ƓL�z ���u��O*i�[-�	~��S��e^����A!O������&���7^�gJY�溕}f+\Y�1�+,�h-Z���������Y_bkZRKt�����_�v�����e�F��Sj-����
���Ñ������]���PJ��i�_���	wg����^��B�V��Rp=�ަ�xK�_������^&#�N�t@d�P�=�M������~|]��q�B�d�����9���ƺ�"A�>y�s���������P[ڠ�lN5�m"�3Ԇ<qp�t���w=a2a ��� �0�ٜ��|�ĘN����
�L�2i��F�����g��t�'�l��$���J~	�%�;�!yW�Q�6F�ʮ�ű�Of
8�A���a4���f1
��;.�P#\�di�~�7��َ�#��{���[
o�4a���NLӛ��Ԣ� ^`�k,6n�����1ۀ�&$����Iƀ6$�}`z�tP��l����y���QJ�w��Z6I0�O���ԩ��
Gc��_'��5���8�%��9A7]�lx�-e+0�Ue��t��Q`Z}��hދ��kGO���@Vd������[ht���P��^*�o�kh��,�x��r
ӡ��{��#�LgNm��R�:��ǘGܝӐ�XxR���ɓ(��9 k,o[�����ZA���JL��7��)�Ҿ)k�O-��e(�DQs�KM��I��$ekY?�ڈJ�{�T���?�{����z��r��F1M!�sz��;sq�<�cw?�[��<
r�$��P���0*�*rC�8�!��C^6�o� ������e����+R��Aڹ���*=��݂����a��?���gk9s?X,R���8�k3񈈽��r�zQ�6��C�ľ�Z����at�l}���)A�-�c#&���5��
a��kW�������v��ƿ��筝+��{��w�]S��q	�#Zc�r�'������4���[��b`��D��Fu�!m־k�������=�B<��������F�[��ވ�]7�Ae����, :ST;"|i�ۺ�,q��W������+�r�3�KigN��I��w�o�A�6�J]=Lu��-]��J U��h�h2�����L�K���^ῥ�'�<�,yY#Jәqxw�����/��%�ʺ@����g�ceG��{���0�H(s&|�,ib�F<�`�Ka�~
��0���r���H�ɞ�3�2�^��W��O��J���&b#7-��|-;�Z@�(�&O�S_�_|Q��c�?W� �����[t�����H����
b�iG�">��~�W9%ǰ��ʏ����1�A�h�oJt͠��_V��75�nX�b�ʑk�x;����&���ݷ�73�~��V��B���Il@j��[���;V��z�m���`/��|���c�x[�)vB�m�w3ש�(�I֠Zd�W��:��Y�,K�~́�Y{R`�p�m���Y�����@����������qd� ����BWdl�hf��Gr�I��*���3�O��[� �qޯX�i cyf�fcU�#���V��(�vY6�`��!u�upo@���BsS�`a�{igSaz^b`���E�c����@��� �0ԅ��T�C��ҋ��U�i�~���)��إY��|}��#��;�<�/�[i�GOnRr�ơ�wTyO��ŸjPt
<e�eP�٬3L��?d��RoJ�rO_{�jadN ��k�E	9a�׏{;53�O@>��9��F ��W���~�aYDza���!�1%�]:��C���e��S��6p/�7�#�M��\������9���RYf���k-�&�ߖw˸*(b������x�|��5���c�_;�6�V _�/��l����+�cZ��S�����X����W�3�n�O�G��zߑ3=n�j;I��x�r\|Y.�g�f�bT7��>T��	9y{e44aIP�N�o9z⇔rX�r�Z?W�88��~{� ��ƏHqm�2�٢�B�!�k����#Ȇs4{�L�+�z�,ε:�`z.K�J��?�;�H�!Ѭ�x$�#޳p�(�^��@a�I0�Q�&�;&��IO��.��̌�Ȫ֧���~���X� jnێ��EI�����+B*�`�z��Ao#x^����"#�
���b�̭�����S!����aPSc�� YM���4�Vm�&�#3���:V�c����"��X�&2<��+��c�§[��W�H����c��Q���Z9��|�:C�t4�L�� ���m�p�82�s��)WD�̘�p�xx����p���W�n�v.�=H�L�מ��$Є �AH��v嵹9�OSz�%�.��>u꧟;,%/d�Y����al+�{{{���9���(t:��kaB:pn"��yN�>\�mEJ����P�� w�5H�7z�4���of88J���čze�LC&+:��~����z�2�	[Թ�B�}YI{�Ǵ����-[��p jb�*\����8�y�mK�#�Wh�Y�RH�<i1�έj�3 rǁ���ǃ�*9ꁡ�$�K�OJ�e�K�Ĳ@q�N:�8jyY���gt�l������g�[����F���s����4�s�ϐ̵e��W�A�㸏�ϿaE�= >.VpYQ��R&M�O�g
r��^+)�7]p�=�|�3�9;���-���G�{ �{7(֔�r};@�h�M���YPo�0������
�K9Y�	9�d�ǁV,�C_����&:S]/g��Sz���k�"ϯ1M�|�	�'R�NZ�"�h����x�������3�����T�6 ;���M>�m�>T$�X�I/�2�I���AGQ�Zpx��J�Q,	�JMnc��~��`e�F�8���)���ڐ	����n�z��}i=���߳�)p��&�G��>��u��o�.s:����d�������9E�� ۡ>]�o䂰@\ԥ��д��q��a�C��+*V����]w�����D�򫆂� �]�nG;�5ahI'
2�@��2(:
���/�c}����Xa�ߏ+��c$�^�z��c�6[��LF�I��Z�8�C���V��P���W��y���~������45�(}��{Rk1�,��#,^"�#���Rx�k�@`�R�!��b�.���Ќ�}Ik�Kl"sD��c �]O,
�\08p��ʁŮdrXh �����x�)6ׯ�m{�{cf���n�ZEh.d�:���HT[�G�F��+�8�ߠ�._�}�����<de�A�b�L-E�H� >�x��?"��_�C�@�(�s_W�W�r�ӻ�?�#��6�i�m�!n���pvϦD|߈1N� e�ę��6Pi��{3׃��~��\2M0'c�#ѽ�J�I0�'By�m�d��h��K��t���d�7:��sk[+Sf���?�d�{�3��X��I�p�A�Eͩ��m3���	4������'���G�'�aN�
�r��/�~d������#���G	��H�IZNy��H
�SQC+���I�ke.�'b�D��X�r�����	M	�+f.gT![��ꃷ^`pA4��d*Z��렶�'����Y���pjK9'�v>%{����"��{����I^$jl��\�,R^I@Z��J�Fڐ:�)G��B6��l��@뜽c6Јe��hL�X��ۧ
񴈢�Kzĵ8y��jT�s��'�:)m�������)��Q��<��?���Y|��:��{����WD$Nd~�l/Y��v�Yl��=���I9K�O>���]}8��h��޴��pO&��H��+}�J�?��~�4{����Bj�*y����_��2So�R�%Ha;��
۠+6+���;�mM�_��5��\`�Fm�r �"�I���f�����B�{�4L>L�U����-8��(r�x����o��4��/Tc�E˹��_�7� �,N ���f���ʴ\��иv�3ǥ^���j�HJ�����N�q(���5&�HՕU��u�?�2�[�>^B��l�Z}�g��zC����;�l�Wp����Ư7����\�����������F�st�m�n��b�\j�]8�D+�nh�O)Oўjv)֮�^��'Q�3&���1gD���0ҧ�#�S��:�Z�7�-��v+7�l�~�r[�w��r�$Y�Ò\h�(`��9�JJBׂ���>��%J0V�x@J±R3��)�5!9���vʹo��l�V�)h���p�n�p�U0Q���j0z!z,No���T��K��H�*w����W�c��5�?k>1��M�0�'4%2KoYJ�tsTh��Bs!}BH��cC�ix7}}JLoG����('/�	�#	rQx`�/�	�
�r d�!�n�"v����P��S_��R�W�����=竨\^�:�+/�g�#.����}�=o��v�|������^s=d��-��$|����>!}�T��/��y�8P �?�|͙\`�frY�FCϮRtH]�*
���Ko��r|\�%4��9ݬ�B����:��Fs����4��҅�=@*e_��� �I�
O�X�,~D���.�X=��x���!+�}��i��͜l���-7`=|�>����V0:;R�$�̬]�������#v�0Q�R �:m����1R��[�)������]6��>J0����9٩�[e���J�,d�g���|V�S������$���~�u��6�~ �CkC��b�Wރ8�[h��z��R!�}[��{D�-32���Etj��>2��ػ#'��K�L,5�nzr�P7
�B���:�CfvT.t.L �C�0�R2�Y �]�V#�9 �	y&�����c�;�]0�#�M�v��=�tJ4������(���)̜�o��2 ��� ���Ȯ����*[xB}^�D�Q����b���o�Һ#�����&��q�Z��kě��R��H�5�n��O���I���q���]�C� �s7IkM����ؘ�Z&+J8.F�/�&�����nr�!�{��l���(���q]��P����{������̅����i�9܄q'��3 )h�/�㜠{�ji���y�+�"=^q��j+�JR�T��5��%�Z_ٜ������������q���Y�f���p�/]��ЮV���hirpϳ@^�plu$/W����&fl�V�L�ޠP�)~�B���w\-����'��M}g�tK�E���]xa���[�sVR���aSꅎ8RF�J-�f
��,)2�"��1ю>˛[icqB
L�'Hr�czۗ��L�������MR��pʼ�{W���2�^�3F�BC���˲q�G��m�07q����hm1D��%�����7r�Lu������Dr��3WzӺ.@��/���8~��B��T�.r�a��6m�l�m�H��ɳpj���±bBt����%��2l�H3:c���  \i��%�KQ�#��at$�z�E(�L�=�N;|Ⱦ)	����U�v�c���XԮ�̶�ɞ��NC�;�(�[�eV	�t6��A7_6겟1Lo���\Z̍iW�Iz�K��2�!'9���J+i��[Hagk���bZF��m("�۫epM�����R�僖�Ġ�*�@Y��D.0��l��YI����l�&"}g���cB�^����]���� 8�����yf �J��żr��E����͚���5��n��(Bj�%s�[:��h�?IyD��KA�bmܖBA�:J�V�@�!�|�ܬ�2IY�s�W��qW�f1-�����������ȳO|(+�FX���z���~Jl�ũ[@UyT��U�������b[1.�<����)���th�
������&܀A� 5%l��҃>��P9ϣ�P,!�ψ����XC�w`\�7ۺ�T�bG�F�Id��i
� ��4gދ|�IK��jYW�ͮMI�;F,��)�������Ta�6o���һi�Q]Z=-�,"���� B�Hd})*��q��.?����:ť Wjw#n�	�@&7�Q���q��D$f
�?o�[D��i��8G"��*U���A��[�WO���1���5T�)�q��Hm�v�+n��(�RNߙQG_��K���ipF9���|Qs���Tꕹ�Ƕͼ��|ډ|���o̔�F�����Ʒ��fj�[KR�G���H�͵�o�V�7�ɧ�M�G���
�V!*�|C.ƻ~A㊧��x��g�t%����O�Z�D뇨�&T�'���X[.�t4����M��^Bp��vj]��W�ɩd��?������A�7giJ!��B.�զlY�O7��-�j�y����c�����vh�/خ����c�ӫP} �ߦ;81�r
�g�ZU�Ps�:~U)�KS}���[F����"S|�Y���ɖ�Oh��� �׬մq�v^{9��KPP&��+�!il���9���U��ƹ(��RG[I)��z9u��(}*F��>y����*ϓ�T㤾������r�뫗��f�:�T�!i�P�N�qDD���h,_$�0��U1��<�[b�"�Y���Eaϯc�zg�*����
�F�����!�:Gv��d���cg,>�6WHH�9h�C��<�K#�x:j+m���w��Q�F��ܤH{���t ~��%�V�hR�������V��%��ZH) �``�t�5LN8�
4Ky�Htl/V 8�ڢU�Ui) xU8M�ѯ���V�����F%�=~29�t��������C��^UP��K֣F�b�ջ�ϧpme&T�A�O,�zY�����)!��v�}ߨ����5*�LЅk�\v���\��E*V�,����5��HH����P��$���=�	�x�Ihr�� ǹ����U��X���X�:�����u�E��39y7Xk���
�a�@az������d�f緧��k���|=��B�����2y��Y�)��\߽�X_w��d�1��t�ŵ��!=�k��5����X���r�8AS�(bas������|p%�C�\3� �(��~3�~��^h�S���YBa���3�œ�9ղ��㵬�/'1�{������M������1+��i��=�r��2�E@T�9 PI��8r��(������R��	�0�3|���X.GL����c��X�"��4�a��g�/�D���ؘ$8l�A_W��Nn�ɇI��큼W�.�p��Қ����	P��>����u/T�`�Lj
^�� ����K>O�&/��T��6�����4U#����F�}P��Sm���d��jI #ܥ�&��{�e�VWGB:2��'�ܹ��q���WD7ƶ}۔I��	Ӌt�X"�=<�>�h���~4!�0�^Ę�M"���x���m���RY�9=
�NVѸ�|
r�I/���x�7�t�����!�&:�|���5��|��,��{���i�0J4���B+VV���〳ޟ�����1�,�F�*��~&��¾��S4�[�.���0�kv\i���9cXͨ�Lt���,�FN�����iQ�vX8-���'(�m%^$����x �گ��Ϗ�~���&���;�)5�Ff>$O%_�T8�;8~��b�VKM]�7�d[tE��=�jb�m�fyHP\6�9����zU���U�Y��wOP��ty�aW�g��5uR,�(�r�yb ���!�#a�~F|[.DY{`L$��ۦ���$�5�����~7�Τ�� h4��� ��ۚP's'�Q6��!��K:��W�C]�7�6뗒��]_�
�(�Jʢ���Ż���)Q�ŷO�,He����Ґ���.M㎁����1�S�:hj�D��2:<z���6��,�[��!׌^�Mɛ��R|�ܳ�sӋ`�9���9��.�_^�-[����Ae!	�]������Fx�S��������-��C�;Bly~駶?�?7�*�w���<"�)#�iF�!A��|=�o`HiGjz5�M�2��\+���m�´p�c���]8��(�"��wp�k� �j|�<�W�m����u.9�C�L`-4����������UkRe=�f7"�P+�c>�������:���k�����P"�z+�P���2��W��0!Pͥ��i�^�_s�Etˑ�k0n)���ۚX��S-���w�����ظ�U9�18sQ�䩒׬?3ި�SP&����#��kdi&(<��v��q�	{�p�3.OQF�;�z�R5T�q�ـ�3�����bP �ٱ5G�vK������y�C/��[E���l��S{J���OJ�k����S�����v.�Un��O� +������U�#�HR��0c.�x���_t�w�k=Փ;�gxP�:|r^���h�]9��h%վBG/�?[�5ε�,�^hUڼy-k�}�]��q��~2%Җ�,�!�1m� ��`l,��0�8[�#����;�� ����gR%_�9�t�nK*�z���Py����^hm�8��k)J<Ͱ��Q�M���B%귗�H�"�!�Z�Y��yrEx [ڱh\%�ٝ�Yb�`�� b������ݦ��yW�Hs2���0�귦!�M�]ד��	/�L��Aܪ�n�G����gL��/1v+��g�N������-tV��>��Z��,] 	��T�tV(�|]�#TQ���&M�1mt��xf���VJ��^��ǉ�b��y�L�7g*ԩeU�T�� ��؎�EG�R6e���2�̴�JI&�j�x��,}�b�������QgɾhKJ��;�=��P��������2��Wȿ�PDw:�b]FDvC���l:�/
������=@IM��!�ŭB�m	��?>n�^��\xe���ǹ}d
ez"R�w�V��p���r��Bֿ��I�L���2~����,R,�Y����b��)Tҗ���'B��Œ��Yzd�F�.��2�L��C�E >����NWzAѲ�$Y��O5n(,/�����ͮ�J�?P�I���1M�ŭ�2�ql)H���Ku�I�< '�ji㟘�����^�<���w����:��
���9���z����Lj1םɊ�#I$O�)"��1�s6&��R�,�#L�o߰��kv�x�MVKl�3gL[���+`mT�V^��$(�\(��d�C�Ý7JP�ʓ�▯2׎m(�v�5#��C;㲻���9��  �r��P92�N��o��6 �?�a\�K=B6�9�'��'�ߌ#|78���F��"��0���՚&JJ�:eN���ET<�),}�P*S�pzX�:�� ��L&#�ʡ�?=��r�.Gv? <�F�&�-{���9�z<Hi�\w��e��Nm����h� �%��
��}�Z�z�%���[~����$��9G��b ��S<����M�N�,0ł��E�ʿ �.�����`��T'Ԋ\K���N��&@�&e#����fm�=��p���zYej�U���� j��`6��ߓ>b���y$��(H��+{��>of�DQ��s8,f�<�D#ۚ�b��ߛ��z�K�64��I�����*8�e���aa�+��+V,��P��U8in��Ik�i'Oa^����H���Rq3X�K�6�w GA�4΋�����{=/�F�]P��Oqg+?���H�:���ه���zO�$���QC�Џڍ��)�u0�#�4�1���e�16�����@l���;����hR>�R�3vQ�~����&�lt�9���>�œA�'�U��U�8�﷫q�?G�0v�-U��#��
_�ϝ�J��~Y8b�e���6B��X�M&~��ͧ��8�\�qF/?'��G���C��c���S����}���M
~Ck`�s��ԍ�@׋�a��W�30!OʭP�[�+��%3����o}���A�	���rW�v�DӴ"eݍA�e;�FsF{t�hD�9w~�Bx�A��Sr~��*`��[��I�b�*����wr�t�E&��9%��a;Uff�n)�*�f�Nm�S����p�،{؊����`�M�Գ'�V$�"g�V�-y�*���6�4������T"���BCY���T�V��5�9P�����Ȭ��q�� ��� ��f���hr��-_㸀�Շ{���<,6��0O��)s�C���w-+Lǣ�$fx6�ޜ\|�W�w�Ǹ T(���,�$;��VfAU7MtY��>j7a�l�1�*�>z��wǾ;n�Z���tR��(�=��bM�-0��Nh�'S�Xq%e���C�#�%��'7?���%�w;x��];�61X���_�&�R0ˠPj�=k���,�	�PGPF�����'��z�mFM��5�@Qh�Iœ�pҚ��^G��Mn-��8�N~�j�GHԷyXQ�1sC� }m���
#(�� ����J�Ձ%��!(ܤ%d!�"�{�p���)O���e)������Py�7��-���� ��%�[�V�Qjd#n.��ͯ�α"ɐ�|#��Y�Jޭ�`�ڿ�tzM>ɸc�!Y:Ckx ;f�3	�ٻ1!���[2M͍�IeCq��&� �gP��F	�|e���e�L�5<oW��P�f�G���[�9G�e�J�%o$ (op�pXj�XrgҫH���_��o=�?����7ڍ�f���)��D�
$®-��zC;\�J�.Ar�p~�����0 �[��γ��IT	�J�{��Zo:/����P�rFUu������4�}O+�A��m&46zc>����a�_c��^G��w�.6՟]���Ql$2kAk	X?ig��j�L֩��BH��	�Y�}=�	��W<DHJ�2���u)
!�}�ao?�D�j�;��K������T�4�8�r���w)�DkIW���F[�YS�D�E�'M���)�m1��	|���zdfQ��r�����B�F��N|�5D��G���=��5�a ��Υ+C����4��4�0�x�ֺA���*�}A��H������-��g�l ᆭ� R��_�T�DV��F1���G7�ZuqsHUbq����[���/XZ��m%���Aǆ{�=�������t�c�i�?��y�`�u|��%i��̯0c��F6��+�ShI��\4[WP�+6��|,g��Xl���Y�7#~:��p)J�&J�a�]e���?)]>Ξ�)nt���>���t*�}eu�R&���Y�rRY����@J?>�C�=�㜑�Y3GN�X1��^�S��آe��ޓ��r(J� ���Qs�5z��I�V��8�K�G:�yko�qx���ک�8]G&?6���y�:�J%x%����0�_�ƶ���z��V�Ԏ�������d@�!���z�4�(�틤?ҷ�:N�
��g/���TZ:�<�U�sN�{u3�L� sN�H5ME�u��n��@�?l�H�_m�އ��P����v��J�G�bj��!eYon\���W���Erf�N�hmP)�U��.wB�+,�-��H(̬�1;�>Yf�����1�tE	rS0ye��~P)a��l��I�%1�q_�/Q�Θ�G���i�w3�'n!_=�1���:CĢ;������,�[��k�|�*ѽ �5>WL�����iT�G^R͑ C
n� ,����SG����Xq�y��ĥ��I��w U�t�@
9AG�T�{��<n7]�@`4D��C	W���WVP7M�����Oͯ�_7Cuv��8�y%vܺ�0�C��Di�w�'�,�ĭ_�GY��ޢ�	�b��,��xD'�x�$� %�2�}XeitB0[�,p �`�uE�f+�{
?PŪ��}|��PV}[-%&+H,^D�D��nA�������]'#Y6�6����x����-��&\���9����_�����E9H���I������Z�9���7Zp�/;�j�_�=��:��*�]�4�?Z��b�tC��#-�[�̃��)��q��/ <��?�A3�!�[��R�o���t�"ОF���7z,+�4G��m�u��9zG���?��0�ޮ���_\��*<3��H���|Y7�2�5مQU�o�Y�q�Պη��`�1��U���{�bJ(f!ya^�u�e���̵r 0�s9m+�uM��?^s�Ⰰ��]�_�Z&,A$�Ȏ���'Zy�	6����3i�ٷZ���)�ڵZ��6���,̼����1y�񭴛�9&��&i=�8�~L�B���2�4%|�S+A����`C�jt�)�h�G"�])u�	�ׂb�FBg��,�ti���_:�Ɓ�C9��

�3�S�l;��\�ca���z �ъ�q> �=.c��46Z�d��lO8����%:����{�bx6ZI(Қ�:���m;�͈n������Ue?V��}R'�����u��GÆ<�[s��,Yy��u��Ο�FQ�?�;P�
4�J�@6.
�Y@�lqѻA���sSK��,�UM����l�4��K��d�*Q	��� �ѬN�c�����S�kf�Wr!X�F�Z�)���<\QϨ,���:����wt����Ҷ���^�8�C�����n���P���d����E�V���T����QW���,�;�Kk���4F�M�����v�#����l����U�Ry���@c�(�*�h5>&
��B{�&F���?�7I]�����5���<P�t�m��_��!��K>��5P cf.[�FO
kczڑ�S�M#� >z������dX=x�C*V�<���`D�W&�_ŵ_�@t���L�/��5�xC�ba������>�p�]6��|rٽ�Lĩ]z#bLtxjs��d��0��.`���������������l����ӯiDD��E��X��o��,��T��;s��,����`Wֲ5ݦ�m�V�� �U�#J��
�2: ~@b�� ���V\�4U�,|�3��54k:j��De܎��2���bSz6��0��^M�9��A�H�� c��5Y�i�^%�6c^�8�[�aV>S����j��18�[A��ق�}B��ˡ�>��	�J����A����10���iGp32RU�	]��,_��������*����`P�鍌��@��i�PjU� e���,]���S����D�I�_r���.'����˹�́yI���4�lY2\TFJ���3:Oi�=8�$��2��3��&PҶ�XZN�g��[��;����@��0e��
k8�)\�@�8�cYЍ��NBf�F��T���ծTU�o�d��G���b	!<�zG��U[�����6#�v�[%Y�w7Z�)�`�uQT[���Q1Fr�Y2T���:���9Xп2B��!A�u���3J���P��p��}��o��0�$8�CXf�'���(!a�c	h1*n�!�;�`����Z��ӊ�H�s�����t�w�g�We�TP��֩:��R�)*�J����S����a���V���D$v�hA�)�&��#��&��{���錶f��õ�e�C*%j�(��-����҅�$8eR)���~�S���Rio��Ef���efEcŹ�D����I-����9h��p�rQ(���co�X$��C��0�t�*(�i��2ҕ�R���p���6���f9�I�i�Kx�=ߦ��:��f�/m�l��D�|K�Y2r������ed� 1�2��Eɏ���a�5����"�~���0�t�=|�oR�}~0
��_Ǡ𡶱h݄R���<I^�H��I�[VW�{��E��V�����6�;��Q�����Ԕ��z�����C\B��{��˕�B�XRD�q~W5@y�m���{�xSl�̹��D̦�1u_F5�Q!�0GjG<�o�����:y�$t�;G�0��^q��d��*T��r���y�s��|3PP��d.�Ѡ]����w�MǞ�cy�g7�g����Hv�\�U;~Ts�J0"]	�5��h|���k6�9uQXg��"@��<�8Zߏa���)`�Ű�4խˈ�m��c�r��0�h^��e��H'��w����c�eb�����"@�6e}Ac�٣�mH�A�t+d}��qd"(/��R���B��O��#
tv*����?������2�ׄgl������D,ږ�˖�j.��Kt��O���4Ą
em�`���[�?t#bK����n֌����L�C��a橴����'q����O���r&����?�2��}՟h!|�0*�����IQA94ٹ��k�o�6,9i�ȕw}��BD��б�x�oז�4��t��I��B���M,wu܂�Ilc~Y��2\9�(5��=�9��x" LH�,*�[���y� I�#H�D�+�S.�u?�m$<�V��8��Ye&��J���:n(�<ln��f�kX�,wGx)�o������bYzV�Ou� ,��s �:MJzI��Q7��FNR�0��(&�`	���v�4�_;��!�롽�HDhȳie�m��B$�h�m�ӌ�SK
ȳ�-S�������?���+�ye���dn.+��3��4_3Bhd�kJ�(�ޞ���+��)�G��0Ƙ7Pɑ[Z�r77�������������dW/k)]y&ff��3�ILf��ևo����Y&7\3G�$���Ӹ��~�ҝ�`O����^�H�wu*�P��pk�x��F
�Ig�L�X$3wk �+��|�0�[�k�����6#>a��u����V��}~�A 0뽬�Ǯ��Ę��*�g_}����^+�c$o��t��r{�G�AQ���Ә�����3������L�p़(��X�c?��cWH�s���U�*e��?�<|My���Q3� ����� �0[d����[g@�1ч�nwV�9ߖ�<Ͳ��=V�c�Oc�1�An�H{U�
H64$a߷���ib�$�7�)D�9 |iy�#�)�dx��c���+1y����;K!�i�7�@�{'�B�~:ɯ��d��,�����`�M;�]Jw��ߺ�iP)d�̤r8���g�c��Lѐ5�X�Ϻ箟��>��ݒ�Y�#H�)��&�q�"'J�j�2�{���g�*"���YD�f���Kt�t��J����
g/���H$���M�7{$���G�{��H�����J�!s ��g�yԠ�sT��$��5J:�4�)hD���-U�b7�`23#39��Pvl|??X,y�}����f.[��4F��Wi�^`��?�~����R1�	'^ͷ�a��Z����Ş<t����c��1���}�yu�t7���ާ��ya�p�sa!��_O�*��n�(�V��䥵�F}�O��Nq��BFq��UW�qd���\�Z�k���z�5��^iV��>ǆUů�߿�\EG�a�V�����ݱ��������.*�&\_*yx�ڋ5��уWɴ��5�r3�7�5k�o��;�[ż��@g�/���1�I�Y�w���b.^��PH�d�E^,��d�� _�8˧4�� ;�qh~SzQ�2ڸjo,Z�=T���q#�J��Hs�SӤ��'i2�{d;�ip8}�29�x�U!��,)��7��7�Bf�nj*�e�qou#�!�w��(��^�+4�^�Ę{)�),���͈��CH���mr�$��X�$�������G`�'���?�̽ˣhb����U���*�"�ѯ-�F�vCA=G �!��I1���'�򠚯)�'�p3=r8��XuN��N1Jq����A�>�"�Gꃲ��Ɉ,M���Ko�ی���%k�W�J5cA^N
Q��^���5�\ٌ�䇽�<�<k��[���Uk�1��^ڗ&��(ǈC���q}��������X�XOj��v�d�R��3da��]LcB�/�q�����{p�> (��7�p�=��x��tJ|͐ыD��+�����^P��f�a7pB��)F���ϕ��	�h�˼���KAѠ��u�q�����x~�L�@�����&��5SW]������C����L��Q���2����[w�I��0<�^	���IrM�sv����$�����U�r�Oa��g�6��x�]����]I��\D� jX$8��_Z	Y�h\�M3pT���I�2G3R��=N��B���l뇢��h1s���Ĕ�,�+v&�3�"�]�l�5��� �a�L�A�DFF˵<�{���5��>w��z8N;Yϊ>|ا��M(�b!>ϧx����B�\Kz�j��0��!6w��*���)�n*��j�۱B�s�9���*��`�q�O�� ���!cH6(0�Hǵ�O׋T��1��ic\�)1��az~	�<�Й���3./���U�Wldǉ��nb��R�>��`H��$��56���S�s���ls�ɢ(��e��� ��Y=��) ����d�P���7��[|�!*A����A$$���Ii V��3U�Za�T��mEv#jeL�?!w���.�U䬙@#��	�}�7[4+�l �%m�E�'�!��/�q�\�g� Ȍ�y��0Ms,_�z\�F�P�x.�m�G���f���eV���=%���Q�
����.�d$_{m�� <�}�V����pr'�If�Ӝ�#�����ж�M]8�=ix����)v��?;tZStx�+w�si`����߹�3<���U��/eLc��B5>�ҏ(��^�e{d��-/�ϘL����pr[�.������-�ٽ��	�}�_�n����{p;��K�h�	��m����RɎ�R,d�� ���?D�$�p��F��i{�A<�C����U|<����5�R<H�U4��E��t�0�-#
��/�8s��<$�^:�)��G���X�l�fTz�/}�E���C6�͓2"���GOlkj�럑и��,�Px�V�hP����������w�o\�zA[o�כ�����=/�?U�g�uƏ��D��]�c�~s��R�*uSvl/�N<ߐw9h� +��n��"�V�e�6S��j.�j߬A��@P��&YJ��Ɏ{��W�[jc�J
� �D���L�%�"1ע�τl�:�i�@��р�w*��쑇cm�`s�2(��e�b�b������X&"qބ'��+�O�g !��\qB3}D�0^Ֆ0�`\�T�[���)�G�^9�p0��[�0�Fm�����X#�OhnO�9 Q]��r�[�g�S2�ˈ7qn�z��l���p��� i����7���Us;�LU�8�\����L�6��0���tl�Cr�Y�����`{�xP$/P��� FHӞ�f9��ߛ��6�Mj&��;Mm0���R�Qہ�� �����O�h��F�&ؾ�y�)ȃ��E{I�0:�tJr��*�2
Ѯ#9!P�Y9V��L�^qȬ=3,ֳ����as��*���e�1����������*����"u���׹�	,L�pzI�[	�J��Fp8"1�a��l@�#b��B_�Ε����[�xJl2/�{�`7x��[��F�Ao�W���������1:���G��A�L�1ꛩ� =����J=���W}�;�@�>�j�ۉRX���qT+�$�2���=v�?)�����WQ���5C箲��-f'�w2��C��6������GO��N�cy�%V�#��+ͻđI������� ���tZ���y��͍�=p�'vGO�%�G��[���f������$�e���7��������~$�"�j��)ȵ���z1��.wn.�?r dW�𭷢%��*��1T3o��k���o���MZb<�!�g
	��yzWAq����=ÕV�PPA�~���c�ob�Z���~fot�;O-�v������K�Z�3�����6��W⸅8mF3Ԅ��a�@¿˹�q/7�f'=�W@X��}�𾉷�ҡ�q�\�Z�-���۱'�(Z� �B�_��ų/��H2�����P��,<����+8�jȄ����r���n"͊��r�נ���%��M.ʀ��`��0��\��~ëT�%N����Umٲ8%�s�Y8ί.#@�F�]ዳh`�iD3��o���ف�ܷ_ȟv�d&\���>�l���4 ��ks�))FJA�y�勑�Z�?��< �j��=��Au����M�C�x����9�c=��r,U��	��\��'է�>��"�RH���%��R�o�w�,	5���θF�ߒ�縒0#��h/���}B��]�J�v�LC&��/��:!�"�_�K��=#����WW'z�蚎�e5��7�E?��ݾ=.��a���陗�9�H�EpT����U�[�d����i�]�fbR҇i�̜�X��ݱ@?�S��Z�:<%��yJ�}��1�ނ'���a��3u�}�����ƆI�C6��?����\�F�ÂӖ��o�vL�~;�{�Zs��-m��v(lC�O7W�DE�r!���겾�l�y��Q�|̱%�D�����o��.���qGi���a,Md?�kAq���#�I;[�Vh^-�� �H��|��[:ϭ	4�Ne��R�y�G�Z�9�n�_v��%w2ڔ�p�ϋ[񖂲mQ_żl�<6I�B?���j��٩ �\)O/���C%`�FU[��5�]�����a�G:��.ZL�r�3�}o[�����0s!�oQv��?��+���o%j���� �0&�kd�RE�*��ئ�:�ָ��=6�E�]��I����1�+�H����jJh}t�2� Lt��u�n6�����_:9���Nd4�C�M2`�/GԐ3t<]5p�­��W�F8j4�t"����n�]��x�����F���ڎa� qYq1��'GUl	ޙ�ꪁ< ���j7U�v�?{�3*�t�*vP]P�,���w �Ce��q6[�'У��Ĩ^��z��h��>�TsT��08ilKD�:X�o�a�oqq�ѐ��Q�!^��fv0b��Bj������>Lf��X�Ӆ�mCj�dd����\ˎ����m2�#%5(��T�E�:}�RTf�a���*�v��e '�G ��-S�`���uP�R��6C6coob������ÒO�z:�O�+���(WzjM��&�E�Rv���PL��f�Fx�]��Y �ݗ�����W,ӊ����i\G�X�!�~�Gu��֚����XبDt�p��5����^�fI/�E2y�<�˻-=ꝵ���3)��aY-0�[*��ґ��b� F61N$������;��t >$@����E����s3�_0��<W�+SM��Q��}�;hhO�����=���;�%�@`xb���y(�+�F2Tb��RL�D3�ޝ�iu_���`�{Z<t�-;%�T|����j6ߔֱ��o%��	��X�I�k��R�q�2����E��Qd��/�����=C7�L��<�mBJ�q<"&J��zˊ�-���/y���)�+�ycL�B���mu���$2�uo6~$��ܤ1n�:L7���?կ�`rD�d��=Z��(�H�e,�ܢ�;):<����?.�ퟀ�����k\�)~�~r/�=R��T��
�,u-tY���7���,i�X���*v��TB.c�k�����Ŏ�ӂ����10?��tL����������tl'H�tQ����m���u�_
O�?��K	j�R�ݘN1�!A#gD�tACe��1���j�?*
B�ύ�9qZ��Ն�5�{(��(f�|jL	B~	0H�����.���T�b6+�֑�lT-�ğ�až�婣ޗ��QF`_bĐ�B��M����Z�H�y,�fR��H~u����X^��S���Â��N��65�w.���~4c�[�x��r�Jv�}F��ZE���O��	���:�@	���A��X)�{1�V�ve��o	C�G� 8u<"������� ��i �DD��:϶�=���N���Í$/�,��p S��]oܑ�-Ш���7����OFv����T�0p�'�U����D��I���_2e��E�%_R���s0#��f�r�VB�Y'�;}i^LIPSk`Cs���b�f?�^�)�d�K�z������& �h�,m����R.���$M�y�\��H����$��A=�T9țoN�Kk���I��~Dkq��� <�[4P�m ��-���u�
R�7�d'N�{u���ە���kC�%��ف!����z�g�Q01;��c�[��Qʣ[�D����>�����
dޏ�:�������>�c���9��cR����P����J�S��gC[6�z;K�d��j{Fs�𒮘U�`�"�O��v�֥����%N��	B�Ƣ�r�#�f��1�{
��{0�E�j͕Q��Žq*��+��}>�x��w�?b ���$����w#L9���4��܄<Ed��*RU����=|��"���3��������_J�HHT��jd"�{���(�ȑ<���������6��	�ݷ۶9�˭NX��I�Tw���(����z>����T25�+�l�,V���l��8�+9Ryc���,Z�ez9O�mV�1�w7J?p��r�\�Y������$�����޺?�b;�bJO���=���}!>lm�3���+h�C\�jy�r����oQw�W�K�p$�F�/	k6�B�n�G���?$бhf�t|x�1�#��y�
��eNh>�\]�"��zl�����e�2�m_2ʙy͜H�dG΃�m�r�"�c�e�APV6b�d�#�2i�W�&5�G��FFTtS���Zl�*[W��X�3rs�)�� �$o��u�����z����;Ifc��\O�3a�?5��
�Y�I�/�g�|�T�_�]*�k�8 2C���$O�������6&��#�{?L=X�'�ot�v��̎��/XqGс<��ؿ�I	�*����rOV����*��Х�3<���M�l诿�,�G]%�R0C����c�`��L�_k�i�V�m����e���s��F��*e�b���V?��Y�39���`5bL��pW���"�7�
~[D,K��*���r=Ò�Y����S��CG��S:�������u�8�|�g��b'^"Ԯ͓�����o�c���m� ���̾ip[@ 7�ve���t F��o�#�}�*���$T%ۯ2�?֎[���m���Ŋd���]ԁ����=��-!"�Ю��{��W`��@�L���m��xo�7�R{���A�˰�ؤ|+����b�x	˷e\�s��c��r��D�VLKz� }(�i�L#1o.�m%�"�����Pec4<�?�⠉8A�x"r|��?��m����������� V#ƐiLޥ�U���MG6Z�����/>�O0ͭ���x2�+�&O�X1��lF���!4���,�PC��q2���*(^2�>Q�D��Ν!v���3N(��
���`����]�p�g
��z\��0��L� �~�J��B�.1C9�C�a���dâ�L2D"o-\ʊ��pC�]k�Q\1��D�YrC6�;Y[�Y��>)�3
����u<I1V��~$��%���kz ���Sp?����L��ٛU���Q	U/���m��G)*�u�)_,�*�x[���w_�����[�N�,Fv=~�j����p����e�jq߇�k9��d�%w#�VP4]�����
���y�W�5p��{j���L��@���r�bV�a�;wp��?�;}�sW��~�K�P�}�$�uH�$�,]f�:�&����X�|I%�"MN�;�:K<��y� x��� �d��K�8&X�7�L�����&+a�������-��.�O�4oe�n�S����npΰ�E9mr���gA��x6N"��gxl���F����l��W"��QX�=����%�@�_��� ��	A���x�a��EZ�I�~�c~����^����c��D�乼�ևr��6�gb�\U3&}�s=`�W´�Հ���3����sO�E��fEf�9��5��!�J`���K!Wn�,+�y҉ց;�����0�U���)�+� �'��EB��℃���突,�Db����5��!�u�~�f.苬G�g-�s���7FfX�!	6~B�O�����R�@�w�#�c��|�:���]���-ټ��z`�S��P����:1��'���P�# �fb�2JƤk�a��H��'�s����h(�r&��c39�#���d���ܽ�j&N0T�[|%�<��T�˲	���G�zԲt��÷J(�},��)B@�g�����{i���9�w�x���㬳[�s���=I@��?�@Ӥ�AL�1RB�qe?8���ή蠇�7�=�G4n�	���&oM#^�W_-�m���^4^vQ��2&�:i\Z"�6��k�cl�&@� iuNM�6��+3*|�:.���`p�����FY�.��Ԓ�PL��t�&�7I�Rძ��rx����k"�$��5�:�u�I�$���Z�(�q=��i�����5G%w�����eD�n����I���Zc|�hn���-���j�!��c|+؄?�����8���.[�UP�e��5�bZ�X8��<��ѭ�`*��h�w%9�j���}��A���7�¹�O�f��?�Dvr<�9�t�ߜ�1L�X�*�c[�7م�W��aG�O��ACN���}��4��Y��A}��8s���ʢ�@��Y�8��7�
�쨴56z2px��?���0�t�D�&o;᰿�kbч���T�4�����m�b[r� Јܝ�~2�F6*�9�'�㪲�
�H�a�..*��_u%L�5Ŏh����pbS"O3�t��a;0���s�����ʹٰOF�(��̛��b)��/+��̅''	�	�D���[�Tx9!,�����l�7L�(kue�=e��ڑ_��2�3��w�%?ݪƫȸ��C!?,Tkq�t͑|d�8��?c��}=�J�r��h�g��|>�U��YޣvK�Õ�@i0'�B�h���<Q�M1�=C)ᨵaʯ;�A����)�"�!Č�&� �T[H�:��;"�)v����n"pҘ ��&~l?M��\mV㡔���*�6,b�OZ� ��J��'�z�H.�$!c_�#(C����=G�U<��~�R������:a�˼!��"G�������I?|ۚ>z%���B/���V:u`��Ģ������� x�Q|�ʰ�uҲ&e
<P��'	E&��LZ�h��%���!��	<���NP�+Poω�$c����d�p����NCF<���U�z�Z!��|�H��3�3D����w{�$V˴\���j�wC��r������@�S	Jg�)���Bx*�ɁIhӱ	��@F������L��*����m5�ԕ��t���Z��N
9��|R����/��ĝ�#��=�ӏ��o�@̏`-hQ6\F(�:X����J}�5`�ʀ��;����":\�#�s; 1ZtS���ݬ[o��yR��2�(� �������IF��Q&��W�$u�,e�`�J�9�/IQ�����t���HV�աiPR���Ƨ�0��ar|�{s3u�W��?�F�W��}T�s��
�����r��*��p�g���&3Z7�\��J�-����@r�-���1���x�^jr/�BL\�0�2,����DHr��ʵ������Q��`�R#��J�ޯ����Y�n�8��ux�*u%�b���/Z)�(Ǌ�wS,	�}^K�g���3&� ��5Լݛx���:k	]z�ap��lR`/Cł������5Z��7��m�w0=�CW�m"���a!,F�,|�=����j=v�&��v�4��R�S�gGp�W�wb�%&d�v�MnM0������z'V��k�\QR���`7�@�E� H�ˌ5+�8Q���O����c�FߠqY��h�2I@���}ַ���j�D�|T���\|}�p8s»�T����۸��	7I��G�cC�������3S(�N�ZD��X�,���n���_G�p��<ON�b�G7l�r�a!�ilU@ryZ_��f���6��U��$��Y4�B�n�\n�e��?DEq ����4�HE4�؉����l���r������)>�u�-`��<���A��c0�k�O)#�q���|���R�}��� ䷹+������o��<��@�y9�&6�����*i��j^Q��0<��U�=r�t�^���$������w@9��X u'ٿ�V#W� �z١�fZd�kF����J�V%������9����G�V��	�!������8`��=�R�alj{���n��р�ag<����Ο%�����;�P�e���1"s��/]X��g]o],+Q��f�C�����QL�ߗ$�8�|SQZ�ďr1hC��[jZظ��>��[-T��|��]�L<s�K��?����ΐw��5g����q�z��J�
|�?��r)�b�!���H�.��]�j��,�&�Rpd�8���@���?oٍ4y{k�Tr����t$
�W6T���h�q�&+�QJ���ԝ��T�@i����Q���ύ�GS�X��)Bn*�M���]����9���V"&"n��(z��T��8!�mX���)HP�3�_Xȹ���d;d��,B:�e��ZO��D���ξ�@���\^�ŏ*����׶����SX�D����U�j4�lI���&�F�������9��*cݲ�J$nR�Ȋd@���y�Yp^ۚ��	mL[�%��L�Ǫm�^F�GD�N�~ �(�Y�yϞ��@�V�=c��_r����u��T7�r�n!ὲB�'�lց?���@���g��ڶ���,f+p�c�{G ���X^-��p_����AQZ�d�.���� ���>�R�tlySt6�@	�Z~�y��5E*��k�&��bo\?��T�$���cU�b�� [ip�?s�k�<�U��gQ��%��OD�D�9�=�A�$v|Q*��F���~�<���b��&�*w��#�N/ѝqM�i��81'�{jRt�0�`�N���E�aİk�#M�ޫ�O<�#5�\�Z��|J]��9K������s�q63_�^ގeU	7p�qpahL�n�&�G[�'��Vw�FK�;��X��#�k?�|7C�Lm���K�_��o}M��m�����ݣy*b��aX�b�Ȩ
e���O�=�S{��O�ȳ�p�$����*�Fo~oz֐ڎl���P���dB�n�g�7Y�н�E�ye������d�q������o���н��� O �鋂���P7��(Ҥg;�:;�k���S��o1�cQV��(�e)�AxDR�4��U�pRM���k`b
5Ӭ/�զ�N��.�����X��<�	a����U�(�۝���{���Ȁ�A3� ��~�:�u���oN�4�7��'N��׬lJ��ښ+����K��T�W�C��<�vM��H�WV0��"3k���)��g����|j�
�d	]8�T������G|�:��/7��lOs���D�h����*�5��8�G8������m���Ӻ�e���)�*Z���q��.���T��Ys���E�Qw>׽yyr �݀�((����$���҄��� ��n��4���A��sG5��1?_i�dt�ۿS dR�P�|�=R�V,ʇ���Y2�qY15����Ѷ�DTX�2�����6F��x�ѹ�����w�曥����y���1�E���HjԣK.��)6����I,��N̵�H뎬w�;���:"��6#?������`I�f\p<����D�\�����r^]���T,��K6`�N����_ۛ�EcU����#��!����I�J��a$��.؃P����Lr^�)�W��ؖ08��ݞ/�pPn�����������P�b���R-,bE����i�������7�D�� �J���Qy�Q���	�G7�]��54�L��*K 1bՃ_t�Q,�WS@������h��VV�|t���=B�b?�}��Q�b{�0�76��S&%wLn֬�8�13O�Ϥ᧳}�o#�(���T�f����0ʦ��uUӯZ_���L��+><�1,3Lc"M��,e�o>f�Ky_�L��T�T�tKP�ݟ���)�%G�@�|jŌQm�\��;\}�v�����s�q�(6:-��-0�SyW��N8�"�/�bt��ڑ!�'�γ�Ͷ��d0뽑B���a�{��%�%��ۥ^����qmp�p'�΂)�O�)�o4�$��ブ���]N�2h��ꜟ0d���q4=B�oV�bcvE@E�dA�[�_t�영�;p!��Ɏ>9�m�4}>��p�pg:��-#5�"��f�t4�y����@r�44�6��%�q3B""N�^��ސ��է�Ϫ�`�RS1[�d
V���f�U��O��FZ����@��.��I~�G�������e��I�-��f���� ��Tߕ��X��\��=�$�p��Ț��+V��O�,�w+��*��̐�g�Vo#�~y�
�66;�����'���&�h��ѧ���[������)ż��A�L#�Cf��E[9���T#�a�wkC �L�Cj����J^=�wN�O��A�;ݔ˶�'���n5��_l�¼(�MN�$���NMD��m_���Y��Au�͘�c$�7xHd�����"]�{�F��� ��}JkdG�; �j/�hk��N�j�T�seGo꼀��w��
�ƍ��qWq��5��� >����W�:�V��ܰƌ���?�Yn�o�nS=^\��*�d1��3?��_���V<���L���~O����������5��c�;z>M�6�e���2��T�L���>L�#���&|��!�Z�W�+�`��+�ծ�a����_��Z�[.5櫻�PR�ag�剿���J�W��ߏo��d��V���7V��"����Rܰ909�[\�r�d�)=�F�=��4�g0�|���) ��-I���ASX?]k��RJ7^�%��L �c����V��Ŭ���ZP�����X�(z!˒��� �oY�_�1U�Q�����ƃ��k�������Ñ@�AѢӣ�'�(숭��z*�G��rm��tA��-lE1���;�FP[l�b�x�D��Ww]O������'1etF�̘e��D��p`|Y	���\��⛫�J7Bv���Z�C��@����6�Pp���}�]�1�� ��P�y��0i��_i� O��E�w����v���(�ZhUd�\�fg
t$�g�
k�W�VL���g>������5-�Q�aޖ�Qh>�?m-Rs�̢S��bZ��Cdڵ^�j����7�koQR�{��in(��Bݓ��-�y�*:��A�َ���E�>���K�PZ$�R*���,��L'`�>g�8
U�6��a|�f�pd���奓9�������sP�������0ۨ9�4���]@L���Ig�ٌ0I�
I��������ˏ:i%�X�u�Bߦ�O��o��{��DM0���RXd���	QR�f|�}�O��/��s_{�J�sC�uM˾6q�9ˣTo.33�l�����E=J�ם4��;�TG�.+���G�K���Լ<o4��w6n8g�>��[���C������$��]����cj��˨�=��i!!k8v%q�����e��"!�B����� M�����$� ��iF����2<R��̬QsҼs����ւ}�=i��!ŏ��RF�����E�|7�zOML�=$ cҀ�G|�+E��-�E/$�:���1~���e*�}R�X:IP���nV[3���/l��$P���mS������G2�F�АL��R}���H�N]t�W$>+||qHy�l�@�bg6G,B6����5o�����8�|��ET[h�2�e�)#���Dv��勋��ώ��eE����=C*
����
`�z|��1�/��s
eU�����n�������.b!]J����W��i˹H7#g�X�Iו�j�Tז��L)P�>��|@*����¼\Ea���@Q>{5���W�m䄅߱�J`�fu:�v��\���e�l��^�$�Y���C�����NK�@8��#.'�Ꞣ�jblK8��B�� �����I�i1R���]�x���,?�ũ�O-k��8������h5�"�!��9�	�s��]�W݆ E@�ѵ�ElO��H'��O��m����ٽ��|\�l�}��xh�r���搉hP
O&ȴ�En�6��كڤ1d�j�um3��r�@Y�������m[�4٨�<d��b�P)m6x������A��/����Nq�m��UJ�銙�t��ӊ (-�٫
��f�{�3��S+���`�9<��4'}��f�Q5���?�t3���DyVg$l�)�ţ
���󆊪��Ռ��WQ�~���%WM����KI���%(-��%\�H��>.�k)�ˇҶ|��	I�j�9Oy�b�]�B��Q$��,ض�G�t���S��[����
�rlx����F�2-[*���R�;?`��q<z>�N���d�hbK���Ha��6�>�@������NUR�aKݖ�� j��Q�ߒ�i�?+��"Ӡ?cXY��c��Q������u
��7��zj\���a���0�K��Y�w4-0b�`cO�%n���nm�#&��nS��u���I������� 06�P����+s"����?��s��<g���w�**�Wpd)q:oG̓�Mw����NN�����Ӭ�Y�Q�4��G�������o�A�n⨰Wᖲɗ@r��A��]��|y�f���:Mu�։��^/�k���'�k�-��j��2\�ki���;����к�����G@0�lݓf�T@Uy���$׃׋��JW����>v.`k��K�mB��2̂	�VR~^��݃ *�"�_e���>�E��h��?�S���>�)D�cB}rX���e }-y4�a�Ĥp��z����>d~B7۩k�	��):���-j.�D	�k���u�GQ8m��l���"�/$�\|�da:ǁ�������v�o���A&�HҬz��Nc�"�����(�m�W hm/?tn��e�.�I�?A��Ʃsx���x���]�Rt�t�v�j�b��Q�$�E��;Op>E��!s$.�Ug�#��V�xE�/z[��<*���
Y(x^3�#����������!L?č_4Đ?�r+�NR��{ټ�.���A��іL�7��g�ݴ�$���*����� ��Ѱ+�rY��Ȼj��:	d�S��`q�Y@fN������� ����Bvyif�3A����#^���������Ľ��C��� 'y@�|i"����# �G3�D�ϏK:���zD��8M����H��:�@�x=����9DN�$��O���x��C�*�x���h���e�{�b�~�t���;�l@
C�N:Zo���L��#1;L~�wlut�&���t�q�	�O[a�u�j x��i�������ܐ�Jl�x��(,4k#��'�0<vAH�\E��(܀ΒU ""\b&�f�A���>�hҔݔ ��5��9MU-�����<��L>ݳ�V܏��\c����a���x�"�`w�Ev��k#"���������z8L/�؅��n��攄Xc�7�n�"q�� ���g�� <>Lk�sc�>�u ��ctA$���P�`���K��s*���d�d`�|�8��Of��¬��L�Qe�%	M�u� ��� �����L��68-�>Z<Z[c�{�5e\��Ng��5�7��j��O�7�)M'����h���p�
B�m��=�R@�pCd��骋��9���ϘەK��P�l9v�"e�\u�.�o�o)OL�[�F�D�_��p �sr��jr >�9K
)�0Ulh��BMz�$Z/�W��Й7�Li��2���3j�l����2h�o��E �^g�dޭ����Q�K���*�+��oM{�+4@�/��7rn��ZO�Ŏڵ��`�NcUԣ��㲒��W�8��;�;ۗX:�7���D��3�tC� �WcG�K���:�9����2�qҷ����>U��r��xPic�����e֕�=�Z�ݜ��K*��	ē���l���i��2m���;�[��{�%V���Yt���J�B������1^��;��1�\��xu=d���M'�1��lK�@��9c>?q���ǩ��v�w.�O�Ck�;����� uce��!����<���u��4��A�o�n��=U�v�R061�ŧ٢�o"�i_��\�r��,j�3���i���H��:.ʥ�}�ed1�Y!s/1�	�x6�]n5_�:I�d[�Յ��FV���h7�nN����*;����u��*������GJ{|��a�3��8��Pr�|�$.X�x>�X4/���=����t�o�&5��M�S��3L�V�j�2���n��W��A|"�K���/���?���O,|���#��T�׆�2�)��&��C�Cb�eb��>R�S�{%�������s�u��)b���i�#�=�ʑ#�'��M	z���n��o��G^�I�:P����F�}��"��V�,w:������⍪հ��.ݫ��m�'�������P��إ�Ϫ�y������dbG����7��+԰��ynx�w� ��_8�o5Qk8;�}��\;��m�Ŷ����<x����"���'֚B�9\0���%�/��f�CսB|�V2�V�Yg7��$Fl�n�e��>9�U̕�tލ�
�|��!Z�Ԁ8�-�Q���	� �^�C�	��2��c۲�4�(ig?��\���tN���&�4!Y�4���81ר �nyˊ[����,���ɛ�51[�w-��aZʻ�\ח����n#�2�u}Fj�5���_D4���,��m��^���'7L��R�UЉ������9s�9B�/�ڥRɶ2n9�Hu����^Y���,
4���/#Z4�N���!"���4�a��>kp��S}ht��8#w5�?�J1i�g��L�5�P�˂o����mԎp�ZNL>:���n��
�����8#@��a��L��k�����3�U`�z�O���& ���r\<�´(����qC~��<���B���80���)k%!R��)�N顷��P�	�q�*��Ls��2����k;�Y����ʯ&�'.��&,�du�r��JAl$��L�S6�����h��X�8�D�Ҳ�4v��.hq*��eRx���C�\�a����9p��
`Tr�;P�#&݉�a�,z�B������+�Bu��Ju�ܺ�i	b��=��y���ﱵը�nWj���%�)��K���G�O��SUI$4"�ϸi9�B;y籤qr���QВC2#�[gA�Ƈ{�1;j]�^�g,{��v���2���A��_��b�4Ġb'g�*\B5Gi��2[,+^���(/eR=�?�Y���
����>����8����κrkܘ���_�c�C{�A-���3�	ÓdmU�Q�\�V.#Ҍ+o&-؁p���-J��������'��pmO,��+���{��w���b 7l{�1��|c״%9��O�̓R���Ԥ���;�h6��F�-0� }�G�hPb�M��~F��EQ�şM~��R�
��IѨ�{�, �{���9�E�V�(�W D�	�k}q�uC��7�
������7��l%=!���i��48�`û%
�?_q��Y?��~�e(}���Z��[l���6�R��2t'��]5��)�4M_?���͖�G`�+��M������`�HFo�~:�UZ�pOd��mi����d�3;�^�4��o�&`�|Χ9�nƶ _ʊ�_1)�V����F�/f�&vT!�ى��Mْ�袅��hp� �+~�oZ�2��F<<�t` ǲ�r�J��zN#�ʒ�g9�v�4P�U3o�pGx���H��@Ц��/�4Ε�����(�[�,��wU���7��莻�
�č_���2����0�t=�a�;m}�:���8�����������2k�s$9}�l�
5���(�S	�0F|VC�j�=+y�yoT��.+�{u���<���l5�(�qӮS�.���@��Vs
��#gL��!aIpbB�<���vA�|�>�zQc9#���x�0>��f�#�ęl�V�-#@�e}$M0;��k����O�=�j�&[�P��g���g�q}Fx]y�'d�"G4�#���|�)kx�n��h���"h����-C��,�����]it����,���=�� v�=��C�Мf�~�\:q+��M��b�}_Y��
�#r��'sYu �
��!��SVH�7��u��t���ݳ��!��||{#����%�5v؀�PTQ�	f��Gm�����&�z;hp��중�1&+�k���NnB^��G��uz%�'>��lE��!�ٞk�f�DeF�"I�M���U��g�OPCm��U�b8���\��uw'��A8 B���_(IY4�>�5��Y���W*МC�z���U��C�%�-qWS��x#9���H� �T31���
J2 pYc�N�c_T}�q� �9��T�"SnX���C��۞+3n�p����e!�_,�����2���,������#H[�'Y8F��	�/Ӳq�uݕ����W��T%8�v�]f�8V���B����,�i�:��/��ޠڦD��Ԁ��v��pG��WA���}5%O�*�n�io�gl<*�S6&q�tkH������^fَ�M��ٰ+C|�'�Un6Ш~��Ƚ�b$?	�g��gMzL����o�Qܐ��_�1��9�5v&���Z�����"=��G��p's�L$���D0���v��
�a���9 Q8SN �D�%ZW�&W5��#w�Էؑ�w�y�ԅ(A��0u6Cd X�R!����fנ���NKq����m4�*�Lt���	&/�~��*^|��u��_��R�+��FP��T�J�f�.�o½�c&��_U ��noa۠Pg��48p��M"�&�;�N@�ܞj���0B��%J�0h�E� ���u���f�,��^��6z�6} �w	
�;J8�_H�ep\5<� D�fu���"θg,�v���x�� ���*:vJp�I�JW��5�/�v^g�7'U��[���4)c�w:؀�\�j��=zK7�M�l~���GVO�k������Ħ�4�3��r}�����2ؒ������1i�l�p����:��b����	Q���k@n���@ye��
��A傸�T����]�7D���n\���"����P-/��
5���p��C�w�g�v�,�Oîk�B[����]&��>m��g"�<�z5�v:j$e��,ʑ+��V
��BQ�
�L���ьw �q�g�YE���Qt'��J5��u\�A�A��_���|���*��̂�-�e���I�R]�!m����'[ ��NB�6G���e����U9犙@4�Y�7�|cʊL	;�&��B̙�@�e���l��=L�lrC*�}{��\�
��yOm�嚹lU��ámP5��֘�R1�c4{��%ʠBͦ�:��W1K?Ţ�(i�JN�c�`����ǷՃ�?jS}B�$X^f���\�)��QV�16ԹB���g�F�+��i>"�N�p�vq����C�pv�0��ŵ�(uߗ�w<�j�] 9��Y�/��[�>P���µQ�yL�^Oy#**���<�a�xS���˽��p �n\�]4���!����9O���}����9��P|&@�ruĔ�sI�DA�Kg��yy�%-�0��#ό���}�CM愥GH�����#}�~�H��'䆭�5;O
x�Q���(�[���.k�p����"/�U�� @Q���%���
��fY�.f���0TڟC/��h��|ؐaH�Ί���.���ڪz\br�VEVPn�b�#��>��+��&v�t(�����P�;!|�����*Z�����QS7�8���p-�j��᭴B��>��H,`n ���&*��dh��r���ל��C�^/�-�q�Z�wdsP�ܚ�%Js8ɷwt�����wQIǴub����IR�'�v�2����r'!��r�0�i�
�#�`��{.0j�61�����e���&G�[�8=7���ESӿs�������8�G�H�W��
���,�lqjs8�M2-tc�G�~���mN��\e�{g*������&��>�p�����Pa�qK�d7�t���U\���	~A�����Iw��@8��vv� 	�S&�g�r�(:�Iie��mέjO�� M�8S$�i��C�����.���>�Դ�[�����p��7�(YN�����V�1�S��Rd��!�i����]z�4X��n�1��H�]f�ר��90x�i��h4��PF��O?�:�vב��-wU��%��hʩ����Ӡ$��AtO�,'ɷ���64X��@ �ݾY�-��N8&���3���~t�>��y��1� �\��~ā ���f��?S�Z�c��{�����-fG�I�"M�e�ڑ7���6[r�K�s� Wr�]��z���f<�����@l�s	�Qc�%�������b���[9a�n6��K�X1n��@�%SS�/�0B�B�\s���=�l�!r��\����G:�gl��_��C�y}�ۣ$�+�;��CHA�8������S�C�E�����=f�S��{!aUvUo K�Vı��&zj�~���`� +N����F�:�����B���"�Y���$�d�2$_D�ESR�EjːA_���X!�٠��A�g�&T�,���	�Y�]�X�3���SQ	:��R:8 ��p�B�9!�3��_G{�A!5�����4N���D{����-�� 5�=)=]ԫ���^ۡ�IH��Χ{���3���}\G��7mm����&̇���z���v�6�����u1}�"��z�(q �x��T�^>��w�l���w-A�����w)k��D�@Fk���/"�9]!Z��2�;���ekU&��lZ`��6�l�;���0C?��=źk�4N��ƹ� �n G����D�roձn��oa�ܽ���-���'�K��u����v�`F�)�����~�l��~��ѭ�4\��#w$������cgo\�<�-[rwǭF��Bp��P�tg����C)�j�d��IX�w�YB�¹�Ʃt,�#�;`�����Fyl��u�w�=�n��2̌�C[��,,YcV��c�E�|<�N���8����x�&j.t�ķe�f],�L�.3/D���)x�O �=ؿ��x��;�cG�u���F�^��N�Q(S�*�net�_�̔'��zg�>�N�C!�2�A���?�gg�c�D��Aاk�P�((���[j��Ofs9��<�k�VRMqU.-p�#C$�AϬ-}�\:��ou��%��-��p3��?�4�-<L�i�eK��
���m��[��%k�p��(z���`�'! [��u�M��uĪ�W�F�e��H*A��Q�S��@�Le�h�3A%
���1���(��Ɉ*2�zK���]�;x�l�S-�FY�Z�c���Ϗ0u�_���a) :*��mF|�� ǐ�����{��"�^��"�*!�!k�uSZn9�ӵ���j�8#�Z��u��ܠ��e�)%��
2��S#�6����R���M6��<�b�H��}}a�t��.b�+р1c-9OgI5�C�k{RȠﱗ7�aP���8����K�KxI�+�E%>%���U�<���>Z�:�,��%S2�; ���G���"��e��%��:�ư�S����*�ÃR�����c��u��~� �4yl��?
)f��&o`\7����Ep��q&t労u�r�`��c�2��K�)�����F٧Cw�7��)X��;�TXe͹�j�hm�1�P���ז�w������;���ۜ�uyy@1REd_���X6͌��jh�#�09���l>�2�	i���+Xb�%%\="��(U�P4n���������ނfJ�D:R����~b�T7x��%�`)T�)6���4�G����`�l��'[�s �TO�G�0'S���J���3�S�:����ٮX��i��$ӏ�7o��Z��1��V��u���@��c����U���8�f��!��B�	�o�ʒ҇��{��ߺ�q�H�j2[|?�dPko1Zg��0�)���ͅ�k�Q�Þ�ݪ����Bp�'�F	ܩ�f�#�-B|;�P��T+�)�a�L��/-1�4q�)t�t~V0���p�/͸j�m�"�;P��r���o���;.��ۨ���j�_�,]���Y����0C+լJđ��~��<�W���`����HmV��F�C�8K�,���c�Jҳ�K�O�n�oF��B�5�3Vs?r�A�
S��w�C���@��C�b 0�6"sh�;�R&K�r�J��v��\��F����2�Ӹ��ʔF�a��~���FlD�mɂI���Cp���D)@p�a�V�(��Ԯ7�ʝ�dy�A�t)�:��{-d>�/�MN��:9nӦͷ�w��h�(#�W�,3��OO��Z �br��s<I�$�J�p:��9�`Y�R��csׇ`�.б\���T����84<�W4�b0D�ۯw��JY)�|����K��^�O�OuH�����܆=�_K	�_�J�ZR�Ա�����¨O"Dl��������ix��d�0�xt�v㤕�2nH�M�!�����#{�g�d�x�H#� �
��D�}j�����%������`���;�a�����,L�O��~Ki�/��`������<24�j�G�W�jG7� ����+��&�%R$T窠������/�R��
6%�C�aS�B��
��,c��h����Lā:���t����O����9%(����,$���)G�O��ֽԈ���J¬_ng�K��%CMjp�$�R쿕�Z��k�Jx�%��!�{S< `��Z��v���pjpέ Sk�;D�A�B<o���q��4��������9�w��05�/�K�vEz�|��`�9=#�7��DM�q �$�dM���&j�� H�����`@>e�}呰c_���?�:
� �|_�X���6EG�+�g�2]�݉
l��ň�Q\�I�Fv����K"J�L"�d5Sjo����W�[������s�{\�f���l%Ȱ1x߲��VK
���%�L� W0EV~���\�E51+���o�e�
�A���U��{2�ٺW[v'o .L�8<?��E���a�A9��C�3�yC��/�C�[ǉ�S�
}��<�O��!�N�9	����.�s��)e3�3�X��n����������ccj���I�T��q}<%D9���E��Y��Fw�����ݔ�;�����C<峤��DFŹ����OgO�}�HP�`� {sc΃��'�S�� %dS�;wg�΢N!����Ph��tc&Ֆ�EW1`/�f�������|��T��sY� �o[}̃��0�'��}��9�
�p��sm^��K]��+�	�o}b�����_�ѭ^�sB�u³� :kR<���| �Ӽ����w���+�J�;K��82;Ct�EƺpFH�+�NN�3���e�/�8;��]ۡ�zB6O$�f_5���a�^�W[�{^O������ϼ	|��3 ����p�6����{�2)����C��=n�f9�fd��ب�@���6�U׷��ӗ��$Rg*Գ���H���g��ʣR�=�&3��9D����$5d�S�dZz�).�A������]C;X��E��7�[y�\磽�E��~d�A,�7_�o�������f�����\�V�K:Gbg��X+X�J$����Tz�Š~(���A��up��� ȵ�ad�M�9)��ۤf���7:I��aŚ��b����ؘ��վY�e5n47�k7|享'Ά��+?3����:�	ց���z���<�Rh�r�8��[��B�y<Ǎ)k��O[Tc�J,�?'���$�䩝J]�6Kusd+��r��Ɖ.闖�Na�^���H����!3EX���xP���z�3(������q`൅k�.F��{�|s,#���D��������6L�|�d�!OA
߹e��rm��BE�Ч߿�
��Y�l��!�۵_�Ojm�G'��,�_�Ї��!�m7���+��F	ҭZ�� �mm���H�y�j�d��+���w}�ޣ/)��{4K�zIA�Q��E�aЭ��-�L�lB:���aP�׉�U�~�E���`���[�9���Y<$n,N�_�5��Bc�/�y�S����U\�������5�0�Ħ��b$�c6����G.P�֔ZG뉪�_�� .Tன��|������ӝ��l6+�P���# +����g$�m�RɋW-�Wم��Q�x
Y��4���Z�)����|�k&���P�z������ۊ�"=�T�*��+�<�eR��I�"�~����h�s�L�W0�;��?��+�˫t�U�~���=Z�<ZO�wWF�fM������.��ѣ�4Im�_�;�Z�e]h�&t�Y�k��z����	�}^
y�p��Ng��|���l�)�v�c-+���n(�NT\��j��|�����+�ݲIR�s�A'Q?���L�9��@Q�ʞ����x�馐iHO�݌A�K�����JeN���t�%1&&;�o����zq\��n��z��r?d���-��5��#!�.�+���ӝ��R����2����G��gū�u�[8�Ɖ�/� <�l,��i�­~INƜ֗/k�xC��}��ʲ�s�Z���>��P'�~Tc[]_���0��S�S��:(�m��U:�ƞ3T� �ׅ���r8f�*p�
C��u;����عS��v������]��� L
!E<�*`?�,]�&Y#J�G[��=ް8��T:�7��-�L�ˌb�?:\�R��Ng�2EG%)���:���d�W�0����Km�&\Һ
*V� �_r�p��)��ov	�v]��<�r��p<���d��O��G;>q�C�x�u�O���XMR����6E��a`T:hRigɨ��#D�]�Bz��RR��ߩ���Qz�v�8N�3���A��*�m���T��/q��IQ�������E]����e�\�*�>uq
���<&<�L-�e.">T D*s��m*Z]�~��K*c�A*��=�t���ǳ�0���Hކ���Is�t�dhq#���6UE"�5�t�^�{J)F?�y�icf�!ݕH���$�*���R��Qcm�,kǔ����_gs=McF=��Y=�������%b��Ն�%OM�=K�i���C �� �[9A^Bay�6�n62F3h&<�����e�gH/M�����C{r��<�%\I;b�&P����Y;�l�GE�[�z?�.f��N�7vm(+h����V;o�yy<���?0Rۨ��v6�.$�T���c�3�jyi��LƎ/�w�$q����d�M������w�^���b
֩����]Ֆ�|Ù�7=g&!�mM�^�T����F�S�_B.'N�q"������z�S�s�p.h�S��z������&��	���W�%i�!��$��xC��]�nM�l��߿�����H�����ǒV���4��iiVp�v����/�i��];mCxI)z|�FAtĒ�V[������>�A�]f��8����1�aJ��>j$L�{Q�1i�#aʼ��A�}(�A~�r�}�6���N��!;�`Y�0�R�:���_�]�JL�g�Ni���A���1sTQ�<����C9��F,� ���u�V������Q�^hԦ-�;�}������'&Ł�p��
�co��B�i�8{��hR�f�,����[�"$-�E�wJkqm1q�Ty!��K�V���d�H����ub*�Gv3D��[&8��=J-�Ԉ�8��[W�\��� w�3�|�CE����ւ�?��Mh����Ϩ����/�Ɨ�G �rY�Mo���U�����S���슂&�\������L��&3��u���p� M�2e���QFѝ��Iܲ.�������o��x+P�|&߯��)�?�����)#�p���(an0ȟrjLhEKҚ9��еʫ>LZ���c�ˡ��jC��V��N�͉���v*���/=�K�].�/��=w��2r���<�Ƶ IJJs��*)��P�Ȧ*�,@�
���r�1؁�2����+#�]����kK��-� ���V�M> ��x<�P�|�t�^	tDp��(ݫ{1o8M���~O{�J���^u�(��ۖ�D20�S�,��Qj�80S��Q9 ��D
1�j���P��@RqZ�l�<L`�р"}���"F�C}ϧ��^B�c����cF߁�;]z���=���R+���is�+����)�˸���:Şz|�Δ�������V0��H��S�R��oX5��Jg�J�uk��v�F���w��(�Ҡ�kJ�(��GK%2�ʷ��9$��D����~��h�hOщy�#���Rs�/�>���ї���s�im5��yNG��G����%ΫM���g�xc"L���8���Z�W�<����5?�
�UO��� ���Xv%��k)���ؤ�����A"nՑ�X�����(��Ӧ,�g�P�:���;8	�_�9�xD,� g�]����/��6Ur����ƿ�-X]yb��7 pp�P8<s;z,ֆ�������c��%=�I��̺�����F���t�5�7�CY_���ޙE 08s��a�9��I]6����oU�����o(���p>� ������U��A�w�g3Is���~Ρ����~؉ۖ��)���[�+MnA��̗nIa��aίd+�%���s�'}��Kď"��!�\f�s=�>�Q�k�i�{�!������8�	_�+�6������%ZJ���]e;4a��VD{)����5�zT0�p�F=Y���r`Ԉ;W�=�"I>F~��h��zc�
]/_<����%�$��.�N-����j�<3}�R�y#�o� `	 K�9���f�0��Җ�Z�a���,O�ky��>b|y׷��� ]p���<������'��f$A�,��7���C�k(o{��d�� �V�_.�sGh�2��x��!�m^�ي����:����,Z�"),��p�����#���	J�<�v�·�q����;��C/,�����砍�j�Z}`�d��t:s $@fT��I��8�C�#�v�Y�!�]9v@��jC9�񄈻��y����_��g�0��Wڶ�d�+�=6�Z�أW��J�-��]6\c�*_o����c������<�`T���mz�U�D�������Ǚ(D���[dS�G*"��0so�MA#k���9~����L���ݞ���1�z���ye㙂j�Gr��wY%��\�V�b��^+TC�M�w�����RI4L��c�1����΃B�.�yp��l��?Fl�_��ˉ�(t7����q�'�K0=-nt�O%�h�J�A�)�j�Bά�w�0�ç�<���S���h�����+�D��[0B�����7�>���sy0ẸVW�L�h��dw�}���S�;5�
���ۏ
k��|z��̟�ʇһ����i�dQyuT�BC|L��?��3&�o��"/�Z�EAd��!�(r5�I��q�j��04K��)W��L��1.��2EYc7���V���A��v΃�k�l�[WN%�vC#{}gUa�݊bb��N�K�u�{(�c��5f��]s2�B��<<��F��Vn~2���Զc��.��)h4�����]���o�Wkz�'��vS.gu&+�'/S��m�:ُxD�1jX�� 0@�y���ez�9�=è�s�0�Q�8!��{�N�e�� �Q��*I~:��w���Tp;�#���Ev��5�
��K�L+�ȤɽY|��^��9"*��>2����W�!�j�?(��5��x��{�5��/� ө̓�p�n�OfG��)$���Ԅ(O�Tu���*�7�%נA������x�+�j���;(�1�iWg��7~Fȃ�I �+��ї�EaL�+��x��?Q���m1�9�|K�@���`�������F�����6�3P��)	����L>5���/�\W�}��ǖSUjK���]k�tNw~�M9������ˈ�sw9�G�<��Q��b����)pֻ��0������
��e{3�6C!��y��Wh�]�AL-h����s�d�����rP�☄c#�;)(t�6�j��eR�t L���?'��0�q�D�6	�-�T�C7ֆ ,4Tkͫ��+m�9��p;k��{
r�Xd�Wa��~�R웣c�W`�s�pgW9��L�	;�ߜ���ϔ��ؒ�X����Љ�	����3�뉯�LC�/��=:8��.���M�*�ߦ�o�	��ۜ�Aa�mf�P`;��lJN�fXxYج�G��u<F�s6~+�ȉ���2L�1��s� $�l9"%��?0*��p
*��XU1�Vվs9��fq�e��A̯�%����B���+���� \��` 5�h��(�k��m�?�3x�W�gD}�o�������B2�t�$�k��O`&��L�*Ld�C���恸�p�7�I�gl�O���Vv_(Վ��P�l*���H�{G������?�`Ԏ���4�΍���hnߪ���?�\���jG��k��K���h���m�s�_9)�Z<���/E
T� RUւ'�����}U�
�ǽ`ܒiXUBƛW6��l�4X�7XU/��_�5�f�@����oqʙ�>&����{g�,�z������0�}���Hv�e���![��X2����b�O"�!����U�`Hx�7�L�{P�^r�R�`���]7_��ublҿ��ϫ]G�(�R�]&�E]��>�[����GvUO6q�x�Iף7��Aw�:�~tg�5�k� �׌�v�k��-LD�Tr=!e�����O���*DV)l1c�c����P�B��/��kI�%�Ijy�%N�h�TH�B:J+n���4�G��"�>!�
S
����s��� W���"�8�/�^
M �����<��sl?���K�m�ګ=[�S��ڙ_)ύ���0WAm�5�$�T����uɝ�Z	��AI=B<=���eT�D��zv�O����B�'g�a��([hhL��,8�����u�b��n�˥㵊R3�r�?O�����SWnA�h�dUn.����v�(�.���]��֜�W��
�b<�ѵ��u|Pk��w����dز+��;)p�X������U�dA����&Cn~�:�+q���Ch8mL-�뒗{�f^�o��}#��*�g���4�9���R����0I�W�{@�E��{�괮����t��$�M(<{���=��$<�ɰ���7u|����;��~D��29��L���O�Aؔ�;Ds�Q	��8�b�QMS���'�`QyC<�k%�,��L1��Cļ��v`���T۰�G����`���9@�⟺�/�9����v*��iT��k�r�v��d�K:��,[�HȒDI��*kH�/��3$^�/�w�	܃���!2���%
,�h��ֈ!�(p׌�o?G-E��y��.��F=��)��7':
�-Ք���yK��2�]�Qu9�6)Q椴0<��9�ע"�FZ�p��2 bR�8���2��Qc�}b(���Z���=f��k������R� �p����ͺ��t�n��)4�6���7i�����;/@���`�Կky)�6>��x�1��\���Kb0�-C)i�g\���3 k$��<���E7(��؜.ayi�zu,���q���/B�L�(eF���jȗ�� �i���[���� �¥�k@�ֱ
�W��h���X�ޏyr?��-Ņ~\�|Ƥ�vDRd`x�ǳ��2�*��В�=ÑF��`H�	
(i�SX@�y��Qă�n�������f[�@G1Mi!�
P�>�A|93�&V6�<���'��0�:x]�uL��fp�Io��d��0B�k��̔�s���_j�1JFB^�X�<ް�/1˧.�Y����Q���@�����E�l]��OiNf��ra�?Xw���o����S�p'�n��lc���mUo���".z+Ƽc���/]�pGڣ���j�!1�3�J|�4����`��w�,��2ۭ5�v	?.��F��F"3�!��~$Rڝ�B]���+�ަ�,�����Ѽ������+��� �wG���F�U��S���)ϡ2�<��@Ɋ�sO�����;�p���ᬻ�,���VbVf��E.�=fa�_���Hcg�l�S��[��U��Υ� �R�������Iူg��Y�^^��+�OZ�����VAvB=�:}_x�7<_��]�ְ��`�;���~�3�x}g"��2*)��>Q�y��Ç=��'�h���@�D徖�#a�˼���v���T� N���y͊E)��JLlt�E�X�-�r��O���{։3��,A�a+O�>��?JhAN�����Lu�yg�5p^��l�H��?BUBi�G��џ�t��J�un{�݅�L�ъd�\r�l�f�G��X����V�#�]�X��d���������ߨ�ϯπ��P�:yX�V��+2��N�H+�g8֞%;�ΦV�9������� ��\��54li�ŕ�Y�%�_;AN��cMAqFB��p�;d��J�?�:�a���B��=TA%�|�a�
�ԁ@fޭJ���x(rBM�ѕ�Sɝz��;��i��*C8h<ɼ�y;4�Fb4,ȫ�.|�u$����BBֽ�o���?��USk�vC	�7��_��L���e�Z�4C{H���\!�S�|-�
��5��`�����Y��X�����뫕�e�~GC� ���	n�樹
������棑�iJ	�(X�~+-3��Vt^
�����x���#�?�W�F/�<��J9������Rnp��Q&��\L`,@�L��!���di%0}c:�A��nFafn�aT�������0�Yֆ�9L'�H����G��	�:>����9�E&G-o#���5���+\��O��w�ɑՄB��*���l3�D���	t����ꧏ��N�V����[Ӎ�k�}����,���?�S���栍uh���c	���=z�/<�4�16�pfj]�|%x����9�����v�z-k8�����4�?�oA�A{`�fN�]I���JTrto��S?�@��/�Ax}e�T�6p���c���#���RZ�������CK�l��.
����I�>�;Q$�'���t�9ӀĔ{cG�k��]�2o�Oe֎�j��q��|Fr� �j� <�2A�@C�_�P�LĻ?f��{�kw�׈ny�+�L��w��f)���AS��|�H�;�
��vN���|8�F�qx����s����_z�+,��<�4c� 2�3����w�9�uN�D��RZz��Qv��7�O�x����Oܫ:������H+�!��ŇK���dCFވ����U���+a�$�'y)�M�j�*~��#�����7Y}�C0� ͛�����rzN�K`�>	V��cB�i�ܨ�;`y!��-���޵N���o(Ų�,��N��!�=H�+���(��8�$:����F�9L~Du7���U�������n�;�}Y��瞈�� �'�V`�D��I���BcͿV�9	��6#]NK?��&�]B1_鵺)�I��L�'���=�	S���� �FARn��:T�-�&�d�oc w`��z���\�;2����qRJ���j��C*�LJ�	F��4#9�^���\$ ��	�-�˨(>El�E��P�`,/�f⮮]H.3�N�⍢����z��c�N�"@}������Bܑ��SkS�lܒ���k�vZ�ۃ���61�"���VՏt���?;�����/F�`�`ۀ�O2&A�͂{��f!겟�C��"qM�i���~��zCW��|nB2h=���d>D���B�����C�I0���qf��3궕"�d�Uż$/F��lm��[="S�j�/��8��YP�2��%6]��;�^8Bs�~�ɯ��ő�n��v i�����M��A�~4#���yч��Ɨ ET��9�쫖�q�A�Za����ϖrD�����ނ����"=\m�,+��u��#�]�l�.�P+�b�ފ	-}&��"XB}�&;�^��4N��D���}E���&u�����"����m��<�oF@�y��a�R����yhO�0y#��sc�K���ʉܓH��'�k\$�?ƕ-��!xA�n?��������260��7z��F��)�� ^�@:�E���)��Jsxtr��& ���rl�k;8^�#[LЭ�^<@�%J��b"�~w��v�X��u�g��#���.�j;��������*�d�w�毋������q�q9��o�P���*���<n��׌eyB_cv���b��۠���arll5V[��gKLB[ZoE�J����-�[��~�Ε��򒫔%�?��ll�zNd��˰n+�|��Bq*�<
)e�|���+����N�i8�L�G�ue���p�O_��^5"#3�;�u3*�AU�ò�$]��t��������F�q�Enu&�'.��(��Y�	t�0����a�X��A�+Z��w�)8�Q��k0������Q�.`�Q
��F�}�ꃥ�{,�6��z�C��D�ոV��ʖJ��,>W�>+%N�z���s�g�n��]��h�,�T�d�3��i'�T�fxB��â0b��>! �,�K4q,x�/�o*�"Ě|A^7��1�u�6�}�o�rS��=�Ia��Xѭ���A>��K;v���T��n���9R�J���<���;�r���37��o�[o��+�/�]�nk�p�b'��7,V��H�peH]FCę���\^���aۍ��������G��0i�c������I O�U��z(;���&�S�ҥ�M{����Xy6�<�^��h�y8����%ukKB-�d^��++XϠF�Mg�]�Ħ&�n>ʏ�9������I��i*dx��G��pM�s��Δ&�8��8#֮Ԛli*u��#)�u�� b��/���:p'��7��
��x�	��I�Y疕���>Ԋ17��īn� ����b�xlN!
K�W�O-k��*#L|25?@��C#.i�H,�sҸK8��u�cDE����B#����^��}`e0WP�"��m�]�,�g���E��Y$��7� 9�Iی#���ga+g��#+o��g���|���7��X*R�a;��/u�	P��a�����m��i�n�-�x����"��TG��M��G��h� !2 Gi{Bn�o���Pm�q)e�X!G����p�>���c�Z'{��j� \���������W<?V^/�2��N�b �{�I�&52eT�W��f�*}\-<���u�\Ȅ����k�r��rlB|rFNz_��'j�V�z��C��E`��՞C�B�K=i��씌"R*1p���g�1]A��5�|�!h� . ���]�^�� ��"�F
m�IR�#Q�"F�����l1߉L�H�G���}׺s?�_�l��G�ȋ�ek��o�B�w�!N:2�a2�{W�&
4�?Π0c����@���G'Lo#�C����M�f�7@:�����	��f��*^�7��ʊ%u��,\�)h�с���y"��NU0�xfV1���uL� �H�ʧ3�2�r�Vj��:_غ�p���&�2�n�^*�'���L�{���v�Y߸͟��2Q��5!鯂�AI4BhD�x����xL%o(�/' w�c�8M��L\�4{.�o�}�d�K�9l�N�RO��c�N��4�߀�����=��w�o#/1����[��hMKmmI���R��)�a�!����]���C����j�񵥵�q���YԎ�Ɖ8U�7o]�n�冣��1z�_�Fqɡ���f5��x�<w���-^X�(��7�����U���>��H��ޒ�v�0�<Eζ�$F��M?��=@G�[ޘ��1=�6�P5���j�lQU�1��$'u��l�:��A�l��|w=��>�hM�RꗺM	=�mg�(1�w/5<��"�1�N1�Dh׷+)��T��c����]�;����d9ٜ��8�Qw\�ʼ��Uy��`R�V���M�s�'�ċ�Ĺ6U�	?���Ց���&�䥙�H�\eC[nu��=�O�jr�[l�r���_�U�#sd��U�vS��/�u�,ILBf�����8o	�Oŏԭ�&���Rnӟ:�qz܄$��<N[G�h5#��P���$w5��P�r�Z`���)�h�	�D�J�C�wn��n|&�l��Cư����oT���W �@�ӥw_���$x��&Ѳ�|��Ek�E��@�qi������_��C&j�?�Aa7�K�k�e�K�_�{:&8}�ϕs�2�z˥�85��L�<JL�p��^;���o���l�a	Da��75�Hn��Ʒ���!xw�L&-YČ/�j-f�`�'{w�����6�/�v{�9=���{�̋:L�f��"&�gr%u��Sp@��oz\=k�����o��g�ٟ��^&�oUYϊJ�b��_nb�;��ϣD�h,Xo�[1RW�4�P���f�E4�Lv|6|D����+/�'����5Oڠ'ӑl�?����6��jt�#�V�y������.�=L��k��k��
�<'���u�^-x�����ԛ� �|(�kԴ<��h^)ϰiL�wȰ 4��Α���a׭��my�ud������z�������ry���K_f"��a����Z��6�!�6=�s�Ӛ���+�`�zP���Nf��(�[�X@�zc����|����s�BGP������(�F�zk�z>�9�gϿL�N񧳞�~c]�\��N�I�+���<� �%�-�A����I���spW9���ψ����Y�Ӵ&�%.m�ex[-~4!�;6�̺7X�Y
�󫵊1z	x�ZԟV����l�\5[�xC!�S�95�wU{n�A�N�������N5��y d�<cdm1�!����A6ѹ��7os��������o�$��s��"u��Ȗ\��]j D��H�#����0�@5���Y+�Y���ry���摽r��`�T���m��>GFۮ�l��"�.���n�`�.}�ڼ�E�Q�HsCj+�Y l6v;��郕g镩������덜9�*M/~���zԞP�dF��
�4��4�o���"��C��D�I��ŲpT��"|�
�UR�$	S�\��p�� �M�ʪ��\�F�^��I�*?�|%ƚ~"4����	@*����uTY��Gk��7/��j�~s�J�Ĝ��)��;-�{�y�<�mL���]c����5��E�jޝ�<%L�!z�;����0>�Je-�"��a==$4WEF&�ى��0���\���^�<���cϫ����,�ձ���6( �EA�������:��~G ��(����7[�ύ��(�{��M�O@�hy�:��Y9/�:3q� ���=��_�l���Uk�|	������W�,O~�9�P�`�ŭ��r�O\#Q�u�� X�f����ć.`�u ��׈��0�T��*��y�]�[����)�U�K��$<m\�x ��a���jR$8LQ�<����( ��Nţ���r\�dRj��X���I�7��\5U?��5��e0�[��?�[BEDJ��e��L��0M�̍�'�x�7��z@�ؤ�'�f#a/L 6���®�p�����F'�!��^57�������LQ~��o�����j�C�p�8�|�[�\w��Np\��w~��k��'k�q%n_+M�5�1ml��V���Vܥ���PM��ƅ?Vd�Lo]R`�Ј�y0O0�@ �X�&Sw��[�#������[���R�h"�s�vS9��j����p}�*f�B�������= #�d	8�$�*�n)?�^�/;ĸ��SbL���%���F�p��9���A"Q,Hs���%��O����X:�P4�����;L8���8��-�D邐�Ž������x3�wK��+��Xa�e����Iq���s�Ξm}�Lm;��{wE�>�i�4�B��fpt�f$�C�ns�"�=7�,��]��Z�I�`�/���(�t/bF����暐a?L�ݽ�O��V(9�G��HӦT��L��P�F�k�|��l��aK�&,'�� `�p#d$�A �'c\�i==���Ѽ<W�	.J��i�X,	]U�Z���Q%p��7^�&`��E�ȇX�����%��	ȚK�v�~G"�y6�Y#�L!8I�ã�q�0k,w�,�a?��C�������z㉞���^>�|F����2�r}g�1e���[���#R���ѭ��l i֔��S��'gd���h���4�kۺ�	�B+��C�f�"�B|��W~�L_�*K�B�N/��?���#��T���o���u���V#F��to����E+�U��m9ڇ� �}ڶ�c#�Z�<W�+K�iZoO2�?��/�F����y�o�/6����j�V�=W���q��Kܳ����Q�ge����cۧ^�H!S.d�z7�w�q��vmWh����Wp[7Io�>��_IZy6��/�!�J_���XsX�O��/Gt����v����(X��L�Uب�`���.���3��h�&�{�"�2e���Y�[�{n.X���W��q8a]��*@:�0Y诹59���EY�����5��J�l��s���hm�v���лR����lم�I�ﭏ����Ɍ��,����ykv!�{�E��'=�Qө��̆�no"���@��F�?E���#Xi�6$��\��S���]��WE��N�N�yr�,	�]���L>�Y$oַ/<��8*I�d��WE 6���7��f�(T�/+g��������塦3�ٿ����C�����f��Ո�����Ok����b���ﭏ��?���M�֯���
kl���.\.l��}�H�0�c�����eL�c�Ԓ��=�<�ݦx^�H�n&n�(ZF��Hb��{xU�t�<u�����t�Kxp�n� ��X�b�!s�on�4wWD8���ylƈ�	� LR���Ă3�2�8(��矀����iYP�_F�Z��wY.�$�^_��X&(��ɚЎp/2�{�[��'��I��ϱ+�8$v���I��e��T��G���1��PTQ�K��T
*c�B~��ז���%�����!_�$��(��p�َ��������I��?d��^���,�׺���M�'�7�QOU����}��q�G_��5N�8A���
��b�6���ݭ�_�y�FS+�����NK�֒��� B���~�0���f��?&�얤Ф��!c�� oY�� ��hJD��zd�A����.�n��BD-LŜ%��� c4֞m�<����`�o���"����ҔeLp�����
����s���(F�p���r�˝���!Sc�!�sp�
YE����I |�'���,�YP5�ׯ�r߱��M:p����Wڣ�߸��|�\9��|V�by�Z�/UN��N����V9�-\�{��:\���6�m�0�5T�߇e#��hJ����@�zk�5�F�Ww'�lI�˖*���[�(�;8p��w|�0��A�m���X`Z���r��vl�߫f�e�o���uͺI� 3��ͣ	�g	�_�L��-�=T��{BX9��� �uQ0�����o��x���&}�<.CD�٧pnK��*�����Nt�}�-k�i�B�-��z��*����(�X!W�G����pHY�=$��)���'w]]t�qr0� ��L%S<gv-J��w�4"�V�Q��?���B#+3��y��\�Vؿ�ݴ�Q�����Wrq�C�h��&dN�BVC���nJY7���ڿ��!m5��b���O�U�*=Β�(O�]���M�~��J�x��Q���&)x8f��{+����s+%�"��7��h	
���u+��Ĵ�y�H��p�e3�Nn�N��/ƾVW�/�~�H�%�i%=5�K��D�������mH凁�;[��U�xl��Q%$��|�&�OVT�q|g�x��sɊ_�!�Pyǹ(��{�����Y,�C���q�#8|�	>�{aTx����N�rY�w�=�����X�f7l��$�ZM8���!�(�����������V���򟹚T�>�����jO25���'"@����9i��`%: XU�igٛ-�H+ia�/�w`�&�S�/�1)���Rhrt�.�����U����dK�죀��(���Ѣ��:�뵂a�zH|��~2��븷4t���V Q���~DV�?�Νcl��Uz�0�qa�I�l�}�����S�C��-v.��)Ǚ2��~U�8�U9t���	��ˢ�r��T�3_�C������糅}�p�#)]ΖU5�NP�ј؞��N�_)Z��y'm4,�(�:$����ŲC(�̎8�f�����2$X0��Mn#�(kю���eE1���o��<��+�H��Ď@/]�V�=(+��	�*929K�{����XG�e��>Hf���T�?��?ғ��-~b״X>5�J{�h*X����4Izv�Ez.�a�N���P{�v��96����v�F\"�aN������>V�2^l�M�>�V�Π����+C�f���\<�IwUM�����νCw2����6K3��D�{˕�L������\�����Eʹ�̓���9�ʛ1���u񯗬*�,��W�]����r�i�9�x٧�N���v�&������������d�^	������$H���=(���D��9�+���,��˫Y�q�h���
��B�a7�#�ގV�/a!��M��w����#g3��a��L������ܳ'#\C���h�-��ꯢ���zZ𨘧.1�I�֡"�b~�IR���UgH_��Z�_,J�'kn���Mq��{i�f��k��DC���L��އ��0bl�;P*�����n3���)��|ʹ�u�2ys!����D���b��Z���>���ქ���1n.G������������ϼ}/ "=� `e�Xzq�*% �J���,�i��&2XDx�WGfo�A�����.��0/���ȴ���\6�զ�֍]�s�yE���b�����F�KvN�$��"�q�c��3Ep7bn�ȷ��� ��p��SMU���g"�r��$:��@n�:N.0;�*^��4Ϊ�>kػ�=a�Y�Ac!��OǷ���v-�t�4�Q�O'��xs�hi��l�N�HerE��n��z��i�؛��C����X7x7�a �لm�x/͡�'������ ��bKߤږ���6�r�xH�iR䐽L�Ƚ��,�Z[b�a�õ�9Ҙ|�T�|�xU�>E�g6ҞEˮ6+'-��X�wdtC�3<�����5P�޲�|�������"9����X�	��	��$������f7�1��r},W.��1L������?5��6i�4&��k��#�����/E�ң.��q��b��E��[jy>��\1�h�D��X��}��Q-���,(t�(�6(˕�3⬮h��G@���7�p��/��p�H�|�o��zl>g!��D�]:[p:;Bo�!�CƄ=��p?�NmЌ�H����L$9[�Ji�t�f�ĸg�v�W�V�M�.UUUrqO �Hu���Xp�Vq�Ӕ���؜I���ɼ���"�d�qߝ��ßɾ�%\G���{��*�L��iw���*|X��3� 7:���
����o��%�βI!�&��9�X�)d��%ި���QY<�N=p��2��G�{~5�;"�Y�6�r$K�Am1�X�ICU5�%��A��j��ބR��4rs]�f���J��1%�t����Ri��>�z��v�NĻ5t8��χ�k�ے)���[P�R�PX��%s����`j�b��ߖ�=E�s�	� ��{�_��M���O������t)��a=����i�g��g]r[������K+�]��s?b`��ΙgL�7�7Ϫ�b���Z2ۨ�Whx�VޱA�����t	�!9�8�ӑӉ!�"�nľ���sv#������?l��] ���K�9���c��`�l f����%iu�$�̕�rgs�������3�0�B�Q�ء�S�lk GD��{�����yz���#k����ki�r-/<�}_
DbV!�`G�@�1�5��ُ�=�W3�8t�m�����O���|��3�}�]�4�e�J��Σ%W=#\�bJ)qZ�%����nT@��"�����_O��'�g�#��|�p*j��c6US�g=��8'Ь���sm���vp��#^�N=;���/���#�p�mGؘ�Md!��=!~Ė]:��B'�I���I����<X� ���u��]/Ȓ_���u}\��\ϾذԾ���8vŏu(h	�*��>86)r��6��h�d�
\�����]T�z�ue�AJ�Jp8\)|!�Z9��v���U�wt˵�"��1�@W�����d:v9��&)e��Iԡ�J@7"m�)�B�<g�S�)��z��Mu� ��6�oP_���������òl<�֗��8��o3�ĬO���b���7jF[�O�TO�A[���ӕ^'+ܞ��gO��%�kk-+���Q*O_��B<C��n�ʽO �LczF�/�T�ʜr�J���1��j,aŤ�!�ukc_�~�4+Kdfj�_M�?a�o>�L�J�r�����σ	@�H�Ӭ����m@Ό� �TgX���A/ټ-J�V�a�$V�B���3^W�\�M?��/��Q�"���N�:���G�H�?������vg��!2�sHWiBŚAUwX7^t���,��gE*3��o}W�̅�=�A�{��m�5}��L���=�h�w�"�"��"2��U)����>�<���C�I���S�IDҎI����T|�_ ~k�K� ���=S>���̄��8��C�ة@����e) r�X�x����/:+�S�����U�a�Uz�-���db��-����9����7�J���������)� v?R�nbl�s���O���>}U�j�XW�>5�}y�fFz���V�A�i��ި��`�E�i�T��z�<�-�����#���<���
X�4A�f��Z)��r6�kēbN�����Y�H��<W6e�G�)���C}�q�9���0	���B���yQ����{)I���L"����4�@W��6�V�\�T�6'ef���r�k����;��_�Y	Pg���T��f�eک�䖈@F�P��MF`
���n�A��A���{-3'�sT�aZ�8�+��WC(�	��=⊻��# �plQ�Y�6=f�ժ����:cSS��lП���
��2���Y'�8���o�E@�^�W�Q183.`����QE0 ����'���D�W�|�$�Z"��@��-o�c�b��K�����0"���R}O;8���Z��A����W��0�!�Q�*�"���)3�n�O���3%`�cҧ�%�v��%i���#��I�sާ���]���n�w���ehc�m���͇���<)�wf:��A�(�5���L�Ы��=�S#Z��������88�^�ݷW�sS����
��*1S6�����f�׮�R|�a��W�����P�g~��O���[�]�V�B�u��J�2缺}I�$�w��BǱwXqc?s.��H��ov���.z޸������'e����Sg��]�13u���~�������\y��F�"����!�zŘ��+T��<Ը�n�4썣�W�rEŸ`��ʃ!�Vi��wAC����Ϸ�8f>�:آ7��u� ��c��N!ݟE)�j����?`�#9ر�������f�U=��A��3�/Z�9��M���i�h���6�c�+��g!�^��/����
�ɕ	+Ĝ>��s ׁ�>��Sg��
�o��f���I\Z�?���#~�׷�E��T�G�CypP�"�s_�'M=g	1����+��AEW'c�㻶됯�Ρ�?2��uO����=C�ј
��wj.U1�������T����}�(]X�[�w�����Q�m�T�j��$��w	���ӆ�pG��!����)�}��C?�����J��q��c����M��6ٰڡ���8L�����=8�z�?I��|�ھ�?��n������M����X�����+�3z�6��hk�y�=o��[v��Q�{H���Y7�=���� �LǓ���J���e�L<j�w��?{"�3��.�B �}��N`��~���fƽz��f���5��S=�؜�U��
���:�����_����q���٨��1M�>�c��W��*'3�j� e2�Qt��a�G Ս�3��v�	��6���>Ĝ��;n�r����bRp��v?��i`X2�G�=T]W}k��l��h��۾�SZd�Vڭ��sny�j�t������$��c�m��k��)��f(�"���(F�,8u1��t'�T �����?�5�s��}*hQ�I�VMMu�	���.�/�P�r��v>��|��*?7��Wwjq�C�f�1Ʒ-�J�V%eq��9q����4���e�����"v����?�$\��=n,��3A�7w0�fT�Ÿ��~s����y�lT>π��+���O���v���wS��˵̾*���ܶ��*��q�5��96��N2F���yZ�j�0U%�Yfxv�)�#�7�%���!zi����C��L~�f��p^���oa!��#�x�,�	��D�~����D��fk���3aLÈ�����ڻy*�pa!Pr�X2���W7��)�P�^�h�Y$ee�l.�Ѓ��`�!�Bk��\�@]e�c$)8!G4U�(����C�[�� �����;�R;X�����G��߻�W1/|�]��װ0��QC��N��Sש�)�(;��Ŭ$�3r�
���eW&K��<�������_ds�ƂN{=ъ�e�b��  �l~�����ۜ�� =�#.�1.�Y���P�"�<Y�{�B��$�ZA��7x�a
�"��}?Խ��[��	��z���D3�[���k�Gd��F[!��oӥb�����$ҹ�����	��S�C���Uw�~kx�����\J�*�v�@��H��&�	�����Ė7�5��q�?��u�.�q9.��Xp��,TT���D�5P�fY�dO��j�I�@^�8�]��6ǂU��y~��½X�������ϣZzW�?,�J��A�ף?9�F�����P:���u�/���s;I�%ouA���+�j�F���oyk���D���+3PV�T3�Ӷ�E&�9S���?�].e��	#�!��&�w'�f�\�l�b��f�D-Q5��I�DT�8�V�H�%������U�<�����rs���r �Ԑ0?n��E�cA�T�:H�N�í��.D��E�p�H��0����ƜOG[��t* �P/�Jj������Wv��$lߣ��b���6(���վV�6]|�=��ّ�kC{_�9�X�;�����r�����k�Y�r���F�kbX�(Cv�sn�:P���O�D�}�s���'[� ��Qᾷ8Ѧ��iR�1�~�8�1���ˣu���#�a�,��~;�*c鮺!۝��R���,E�g+��=�4P���I����3Q���59��L��m�k�)r	f���\_@7+a.<_�u��U�� ����񅴱�������;R�J�����"0�'0������x�j�K���Z��b0�G�~Eٸ_���	���t5@x�+A���\�C���"{�%���wQ�����9��G�~��r�@`nvtz�� ������{y��A����Z1=XXR�?[^�3�Òn�7���ʮy�	c�}�%�d�H��"�7$E�頦	TV��.��K$��Iu3LC@�z�b6�T2Y�,�Э�^�`��h�C����hݺD@�S[��̄��
���;��q���[��g[k�̴b�/��!�1�����N*��̱J�̒���sIA��:+V�}o��L���M�w�΃<p���-�%ߒ�i'�����j�޾C��<���C�D�M�''���P��G��˫�F8����  ��I��G }��ye	B�݉-���$Gj�Cr�\xs�ur;���3�O z}6�H��ys��.��lLH�'�p�yrX�>Hi�m����������}�#�:�Щ�z�ϔi��UI�]���W®'1ꂑ}ʭju�̨Z�Hȫ��)89�	D~�6���s(�㤣(V<q��{�A՚pX2�'jF�2�8mp�����+;ms �
������}�z��{S�ͩJ�࣢�/����9�� ���
�\���EB7K9���߻����� `d��B��aZ��+����VR���E����4��N�mư���X7�Gи���o7b�C��H/S���&��=]�#�	��"�{;��Zc@�O���b���i�%	> ?= 4��u��ǿ��St[�Q!+��g��܇�3`ܙ_�+6f��{��
`�G�`%Pd`n�s��і��?�n�N���2���	}~��{Ƌ��$�z�K̊Xo�$�ӑ;����=��y+�^�g�6v�VE�.17��W�����&st{�k�a�%��e_hj���yae��NHx��꒒ܲ�Y�(��+�ٛc��:|<���@8jU��}�(u�"b/���l	|���K(�i�t��p���1%#>��֎aH�Y��ۏ��jBWu���y	g3���q�$��<����\�M�a�>�|{��x�=�%)�6��Q~i���4n�����m�]>��@C�-w��e�j�im�j��xwc�Ç��Tvn줣�xc��[��lu�����1v�x&��$�k�V��������	��d
g�5�] h�/�����klzM~�z5Qѯ��HǑ�,�+��}%�q]�dP�"��H]/�o�ɪ$tb��?���RE$�7�Ac����:�'�2�~r|S��9��1	s�,��$ВFr��)�%�{~�Pr���;��H\�E�a�Aho���M�Ȳ&���.*V�. S]�=�Nwe�����o!��ٽڠ����c^�~oУ��u��ɴ�E� ��`LZC�W�V:����cS���%.���t�E�,*I��1�\hmw�X�|�m{�K]��%M#TѐTFHb�����ڂ�yq�u�>����D�U��e�#a�hl��n�vJ~�K�$���.*9O��l��o�!��x��;�:�Ob{��\'�Tx�u�񅁏c��&�|���Fw-�/t��1�D�d�����"?x�M
 2/��m�׉l�3'�.�i�G�R�6����������;!��ʺ��n�:a��6�W�'���<v�1�~ ��o���Vj��ڛ���c�DH<u�%�$8f�4��(
�vS�P����:���M��#ٞ��P=��Ƃ�]e�_p�L�v����q6���1%b��0ZF��l?�VƦ������e�!��{?y�-�7��x�e�~�.�q.��7.���ڢev�:@+6�v��Z}��#����yH����e��H��M���#4f��aj_е^�r�:�dN;��A6����D��rB~������{7��� �s�aah��Vl���I��K�~���'�H>"|"���$�U��{~�4�PI1[�I����
tm�:���g�jX�cyMv]/��:�;2p�
�� }��	���a�_T@Br;�o�[�zF�r���p̡�a]]؛C���<� P���^���i"�]�`��'��3����/�'z���p
�A2JAM���6T��*�;�|�H�S��]c#m �N�k�đ�f��Y`�d2�B���s��\?=�/]��r2I�S�Y�ݦ����،�z�{ cI.�%�DL��hҿ��8ĝ�7�jϕ��6�Sѵ�c������/ټ\�kXG]c����̀���r�O*R�,�2k�ƞ/��$)IVh1�[��=���U�A\䴉wY0s����(5Ϡ-Th�%&��Y��Sx�r�FkF��ͪA����������E�|D�}�D�7U�w�s|?^'}�k-�Ϸ�}ŏO�+�$'�.�Z�C��R�����Ն7Z�"U��o�b��_��x�gf��ύ!�0�� T�m���۠P+�w�q�_��}��H�X�p�<����rj����9��2��=��"��)h��&hٶ$�&����t����M?��!�{��\z�J�<�2>[+�D�lo3G{t���~�mX�V�1̷s��*M��I�,Z�����u�3��嵗.���wvۂ����D�S��C�(�t�/Tj8���<�ґ� �K�Ӗ'ռw��};�ӽ&+�2��2�?w��+�3T#�_��ƫZ����e���o��C#�t���NA��!&Ѷ���{ʈJ�/;[@�4`��og �� 	0¶X���f
��uyHA&w�m�}��$|οc���C:�Xm�Q�Ýk j<�Җ~�	����_p�޷M@�w1ͮ�N�t���9[{,cϑ�i�8�Iȧ,|Ty�Z��dlt#��{�"�0OÇ���)y𔤼�����]c�Y�׷Nl�/�L�!���Z�fʓ�[���^j�B#���oA���&�ϡ>�9ސ[�5�Y�1��^�|���g��VS��-����jZ��Y'G �'�!�>{�5෎z�W�t��[�t�a�P[�BE@�irI�?����3�B���$s���~�I,\6��Oፆ�H�`�2��Y}5-xY��'׈��f0V�>ƈ�G$k��E�����u��LĲ+Ww�����S�a�����>pB�r���P�ʜ^-���C��C����B&�҆�NWY� �9=��V�]�yh'0��zNvxϷJ��TpEG��ׁ����gmK���tjÍ^�����]�]�g����ޟoyf�A��&(S�y��y��F�R��7�'�	�Q:8ƅ������h�oP���>)mq�?Y+zN�U���I<���8T
�	�X�o�+�Cbn���u\Pbז����W10- nNb��¸�$0�)�L��{���R���D�J/hA�d���v�>ߐ��~= �$.̹�IՑ��0���!�Y�aD��g.��k�ynh�)��r�<�V2AGD�b���t�}+SI�}�&ڱ,�=-�?븫�����Z�s=��c�����'��[	�vl����#!����B�i6D���F�=���G�&;H�;�~�P�g���{��<� �e(��jl,�8�諸	�U�$eT���MڠG�wZ�z�5d�]��}���cI�˚����2X"ͣ��
�o=%�壡�H���c���S��Zf�v����"ӌ,l@��3=$�V�dU�R�2	Na�K�+cX�� v_ɴ�6�n	�7Nt%��{ȟo*x��a����!�7����		���~\���B��͔(�n�8�l{���.���-O>)4-�~�x�8{����u����6�= V�zr 0>�x'�g���..���v���/��_@F��M��U���!?LV�b�~���1c�?�*�Y�p�F�>S���h�'�R�k0l��*$:(a!��>�f���I�k��@�7�FD��D��l�q8�s�,4���,�\�L���yJD��?�����P��TX���G��G�;�{������#ѧ�(����u�p#,�u-9�C�
L��~{x��F��M���,/L���l}�2�@�XIXoB�Ï�������X;`g�r;�-��7�١��
g:���pm�s<��'���Nw����V4����1�PV7�;½��yуu\L�w��\Z[ƨd�����k�0N�ė����5b�Ћ�(�>��5J�TsK�*�>\�|����;�7
����PA�w�5�j�8�.�2�Ģ�ʙFؐ�j���	"ξ��lJ�}y��Є��9b�u���:����<X�z��A�'�zGS9X1|!�{\Q��1sĐ&l�qO��<�g�k歿���8���4�\Ȟ~7� �>�.�_�,��J4+�0H!e�����d�#�����!^~4�jI=Z��!�b�?(k���~�j�I>�g^����]�ku��-�x��6�o��I!��z]��S�K�5�DgA���m�`���D��@@c��>Z[$��f国c�7�h��Yަݑe%�;��dRf�&��/)�[�͠FoFP��34s˸�&��`�fO�Kk�ܶ�ʐ��M�Q�ϲ1۩`�n(j�9����S��'���vb���ȱ��=��_��shm�>./H��Q���y�W�~�_�#�4����n8�����p���%��9�*r[�W�2��	X�8��b���uO�h}NO�L�D
�S2Q�I�t�{-V��!:�.�֛�Q?\h��=�����8�[��S#��jji�ZE���H4T��?V�GDa~fT����s�dW���+!,����˗;�R�0�!)k��g��yr��(����=DHa��3��y)�zB^���˽  g���l�e�׃���Z|�n+��I�-��N�%}��i:�nYi�CC���Z0�)�������#�]�	�u$�$�O̄6��]��>��[�d�{�cw���� ����3\�q]�M��@0i��$f8�ٜe�<���$#���o#�ؘ�f��ylٔ�X��k�^:Ry�<���'�����L;�5�)`���ď���������J��.Y�^����S)�V��+��aW�=%><��,;&t&F�RhEM�����7G	^����j|�a�mF��|��lԇ�+���z�i8!��}PCf=- �8Ǯ�R3D���&� S
��;�����S�M'�Q�ҁJ�IA7�Z�`��[�hMMŦN'%�'֓���|�j�l�K���2��c4���5�r�����l%	��XQ03�ܵߪ�-�.J-���<�'�KwG]�����e��V@�bJ^���V��j�I/[���ܲ��>�E$���7�$���z�4��&�N�p؉G�Gd��A��'p�Q6�5^���7 �=^�z3G���*�*�K�G�p2�i�f�Nw2n��#�����4��S�u]_��4��E 7WYp3�'Ǥ�?VN�����Q�W�oOA�*������
�� ��'�яGD��4ɢ�K	9�j��3w���P��,����X�)e��/�X�;��`�A%��5� MhZ�H��H�`�X�ܗ�M��Ɓ3�'�8a�*WL҉��Isa�k�ZfXef�HS�)�6���/OC��m\.��?�C�S0� ���tZ3c\��|�Y�CE����j�9�L��X����p)�.<5��D��f@�.�-��-{���Z0mF���e���|��`��e�é�ʳ���zDh��7FY�,j<y���n�x*��rZǃ�W��c���E�pF��6����q�u�*Vq��	����1��r��g/0�X�#w�P�x �_> =K�{A������ګ�S'1E�m ��e�G��w_ !��m�-�Zߜ&�*3<�F�V�}j<��#Y>��<�U:P���E�`܂�m��k�<� C�6�O8�z-`I�y/�I�6>�F����Kd�9��x��ڒ����uqL>I_����E����n��������1�.��~S����r�jlh%��� �G4*��>A+!_�HX;_��
�u[E����YD����kKGd�7i����sA����������K6��t�^���N�27�Ϟhg����b�$]��jj��-�E�\�����w�����	n_���ȷx��ѷ%wTO>A2Z��/]$@�o= ��i��4E��c�	����끘sP��Ʀ �)J5r%�L�߈�9ZHg�V���o�_H]�@V�W�Q��+7A|�����%�/ m��k>�I�𽟦 �z��H/�g
ԊoM݆D�	���U�NA7��!\4�O!{�g�c��>�	�멉�w�·U��S	���J|��~���+m�5�M�k/�Q���;��<��,ޛg-���v��=����CL�_����
D�;JHk���'�@+_��к�`�Z���|L{���}J�$8z��I�(qE�hk���6�v�W^`��%��9i��]���㍂���,W�VPA8��-45{bJY#����X�=`�}�|[�P9�$��ޡ��x( )��K�J����tL�� �ڋQ�eY�sYL7n��[;�׍n�'4� U�#.���W.�`'�[�}�|3�y�RH�v�Gvq;R<�f���4A�tc�%�1~aƆ,H\e�����;�}�-F[�U��$�����`��z��&�KR�QQ�w?��X�G�UUs�*�#�����^�A��S���Дg�Ch�p޵~[�X�8�'qq�Ҙ��/��Q�LK�d����hxV�"<�c�~2c</IP"�����i$�i��`tOS6�qZF*��m��+�y_��т(� ��W��z9���\#	�x��vh=!�@� o`١��#��>�y��� �CP|�g{�9�v�ҿyMTC�Y�n�t��R�T?���rs����?U�ℎu���~%��5��~!�`d��Ž����3o�;�s���K�#�Kmo���^�!�DH`��R;[� 4�|�py�N�/��/�����g�^V���-�Y�,�~�Ei<L���L�`U#d�i�ͣLG�z��gÝ��R0�T�Q�1Kdw~r¤��!U<#�zBx�=q���A����8,8�"�g+,Z_*"N�)�d�_0��Fse��I9�9�nG�b&�ޠMsSÙTC�ʘ�{��!Q�u2��-lS�s�q��Ƴ;���0gV�ܤ���Q�-��m����A��}�c�l���[b��K�dT�'%�y|t� T��n�VJ�|�sA��y,G��ȢL/�+��p�|t�k�o�4*�~���j˚t� ��`�{��5�d̨��N�~�#��;��o">3;�;�`$jq�~S/�v7,?rƲg��[��r#8,���9m�k7
��*LQ��%6���vx�u�O���9F;��y�.�J��J���83ܾ6��r:Q�t�FXb�ٖ�t)T�qD��)L[@A�t�
?	�M��;i�@
�h�oF�-V����	4��J�������g+>�	���V�:R^ʧ�j�J��6��8e���o,���fK�o�uU������N�u�!�:���$�e�ǎݖq�]N��������1�S)DH�L�1?�p�Sg���m�ϊ��&����J:Ǩ�z��-�[;n���D�
�fe��<��m���#x� ���q��Mt�0��y0LI�cI ���".y:���s��:խ��k�7m:�_?���F�Ɣ��o`H�TQ m�ъ��ȸMNKz:�bk�򵵈�6�'�Y�g�!�g���a����x�F���
�)�����F����qR�7�4�Z���6ԉ/¢\�؛ymH[���QW�r�\?t��)����Y�l�W�%s90��"9���e�n� �e��X�z����6���K����&�ˀ���.��ld�l?�rh��q90���P.�jQ `�G3�q�G�A������J/k�����C	f��&����x89<2��z�SS�<��y_��Cq_\�|�2��%�W�ÐqEzI��3��P�+\����[.T;�1�1ͧ1Y��Z(�K�/���(}y��2Cf���Ŷ�*�䇳{S��O�{eQ�7�.5 ���>%���@{����f�;i�X�΃�Ţ��[�����õ�r�f������3E�5j���g�Ӂ]i��b�`9��4�?�aǸz��W�4��y�r�<s�tI25[sO,YŞ����;$�t35K���F�"mǇ�΄�`�ty��B�lޕ���a�W�X���9l�s�ŧs���n���:F'i��t6R����%֡5w�K��XU(4?��ꈙ�NH�j���A�Z��Re��kZ�L�#vC� �Y/[�o�ܪ�u���}�=^F=�Z��.����_l� ��>G�C9�jRv�h�L����#��9��%"�U�}o�H��v�6ql��x��ҕD�Z|R���ch�2���C(�SB��ݔfOֳq���	Uܢk�D��s�|�X��6��-���R������Y�0��,���rt8o��~Z��8�P�II�X�<B�Ӌ�Iq��	�ߏ�0����|�p=Ns�]��4�앚T,�#���0p;���R�	C��F�yy�Յ�����y��o�"9���Jp��\�y%�G��5�OEK?�+	1p�md�ࣝ_�M+}>7�"�!D08v	

���j�{@��Z��TK�i;�W��Э�@{�z5a���2����'�n�t���Y��re����/�:�����q�!�5���}>5t����w��%=A�n�ɭa���}tM�?�)y����m-/{�s�S��C�@w��5�N�`v5�U+��Žy�cq8�n�I|G54�L!�>p���]q��� М���Oo�>H�R��N�"���������S>b�?�_��X:�"�[�(hk�!$�*Ɨ�{E���IM"�.�^ʓ�5��M�c]�gXP�cWv< 褿��g��P�N��RHF��4�D�!_�]:3 �x�/
o��u��п�-�ꃓp�`/Dٔ�I�[fO��p�w]�b����Xz�Y�Zs��x3�7�4��͓�� ҳ$�3���G�V���[��cU���l��L>��F���At�{j���rc�"x��;��U�:��_�	�/쬟.p�/�vN���y_qxN�I����y.�̛������w`�S)4�%ճ�	-�Q�j��<"��?~�Ow�mn~����l��( ����i�OA4&�`�%W��_=@����2�W#"K¥��t�%��:���	����*}��|�<����v.�
��L�2g��t~/��)-�.(�Ku�~���&�|KO	6�.�~ /�|��=/�;Zʲ���0�m���m�-Dy�<���r��^ـr������� ��s��������߁�v�4��@]�q୲�O�mTmh>�9�FB�]�[�5S^fѝb�NX>0�V����`��ҋ���0&�v�p�tO�~|��2GX�I5&�{�?��BQ�\J�A��LgOf�ߋ��4�l�$J'	�DG��%��S>�XG[��7q�,����
��t*%�]$
f$��Ge���':IO���=��2@�G���P�x���۷4���$�W�Mڞ�!�d��
4�M�o!������[����&��T����u���R��B\������W�r�F���D]��z�����7������K��*����w?�.�;qjY�^��t]r�a&��T-��8	.j�s 0mx� ���0!�j���D���SM��%��ظ�Oh��(w��MI<��)�g��t�|�2�� 6��)��F��P��K���@P�ȏ��W����WCG����j�+�kr�@�ȋ2cJ� �ޗ=�4hj��>R���͏g��� �g�C�^GQ�F=���f����Һ�b�k���pkG�B�"Yև{:����T�ԕ"�)y�<[2���e����Nc���r��S��8��2����������~�����\2��`ߌ�e9vKFv�,e$�)+��D��h*�X$��S-�p:�&�Ņ�i@ֵ�B@�� �(��̜x���9���9���$�I	�~G�VJ�{D�;!��d��<�zְf�¥�R��Sm11d��i��1B��3/�����=й�mDРBJe��~���a^�n�
��	Ԅ��)�[��\dGj����"��i ����
 ������x蠫���x��~|S.D�Y���V�c���8��̳�w�H��6��Nj�9i�?��`��!|��B䓱�犑��;H!1����1ʷq-G��nw̥���(�l��4,���NF�`I.�<�tL-�C�QP����� ��A'�h����-[�&,�RX���N9��!G[J�w���כ�k����ʕ�.�\�I��ky����J��W��m�ǋ=�;0p�':e�@U=��׼"�1쓡Ƕ"/��5��)��[k	���W�]��ߩ_��=!R��n�g��_�YL�j]z���X�~;�����\���W�?��du�y��w�����̕V��3�d�Q?w\zWp�� �{��"J��:�EdY'&�D�
ʴU�4�A �j-�l_b���Ѫp{=��<�|�ٳ}��TN#� -\b���hٸ�$�N� ��s������x
�����ŤG�% �g%UA�S<?��.�=��{Y�*���߫ߤ�&�����3y��q w�P��	ȉ��1�̼����C�!���)�����*�`�<�/������7g_7���K��Uzx����c��-ؚ>���aGTp��Z갃޴��䷌�@,�G�)����$�������{}��E�� ��V�Sၵ9w�ő2f(nX���+{�8���<p'��H=Х��1���n ��P�=�%H���Oi��!����X��&�/F~]�I��ʻv�w��m,�R|�+���
��΀󎵜��8��M����17��I�Z�*Џ�E��p�ѺM��j|9ͨ��.&�-�@�j�m�,s3��5��d�=�K4@�g��h�^O�-���H�T�`V��T���;�beU�"�gvC?���'R%qQb����s�|��`���6�'����jB/���}Fbsā5��D���G�z�`�98�n���/�������u��Dm���x�$��'������+,],�B�r�v��=U5�j��J���{C
��JM�Yi�2]��{K���1(�	�n&
��$���B�,l)�����}���ӆ��ɥ�+4����25E6��|�,����pKk��@���%P��`�$�$H܌�Ѻ� �Oʹ��꿦�`��o�)�d��mR�+s�,	� ��U�X,����5���"�Q�O{�\P�4ȕj���U'@�e���G%*(�w�� pG0!M�C5DR$�fW�^���Y�}�T-�0HM�p�:R_��	���k��y�Z� �i�u]b�y�P#VQ�Qf�.����H����9�2R���������z�r����|���fKor��@�wh��P����~�3�g��u����+�Mh�`o�ڤ/Y�%X�G���|�t�\��Mj�mϪaXB�ݴ��Zg��+�Z:�a��Z�k]Tx���2�_��W���G�k�řH�(ck�Ny2C���f4�/�]�T���Q	��HJ�j1h���~���U�A���aU��?t�,������/9\ �m�?���[��U���`��=��V���E���!8o�9Yw����=���#��7��d1 �'1{&�ϸ1H���`��=꽦whN0s?K��,QUS�h�ڄT�|g	�I�� �I�א��G	��ꮴ�����@윩��A�BY�H� �l��B�/;B{7�hkL&����H��yY N�0}����a�C������\�g��T�I������J����{�'J�F�0̵�B*��"=��*Dp�ױg+UHڐ��ZO��9��][)#(�@y�Rx�a<�s]~Cr8X�	��_)� 0c����[�����V�fl�]s�l���X 4���zX���N����駯�}0�����=n��Q�胭j��z�`x�}ό�Z�ZŮ�/�`����\��g��A?̤F��8���ax:zժ����U3�M��*�ݒЈ��kS�Ź<�s�F8���A���F�9'�՞�j\����nrQ�\mI6�����z�tǽ@�i���]So���6r�_��S�fZ
��f���>���>��\E�S�|��\��X��L8�^��PV�y1�Zr�!�3=yŉ�E�������|�Я�Q �z�>a��_���m�`���d �F6|u�̚���W�sLt8Ð9�qv���m��FEW�Hq��Є1/��K����G6o��Kz"�xL.�N8������k&��Nz���}�t���Ź�N�������SPV��#�>�6�����4a^o�����|i�AT�~E��a+~r�2�Y�U'�9L&�3�i�8G���}�+C��;��rCA��XZ[�m��͏)ΔH���#�%��6~1:�^9�B�0˭H�� pq=R��t	b��B�ޒ�g	����Lk�N&�ت��}�k`c��	?RA�v��| �$�~6�Jv�0]c��@�[m8��3߆�D���;�77j��ob�K��y��F�u�����/SnWH�K�Į��z��V��G�뎪�����!hf��LP�0W&�?����o��v��j)8�z+sN��Jx�p=0>(���c��$�:�d<Զ�n>�>B:N�Rb�9 ���,U�"u��?4M_���W�%�2�Bm#�0j��v�3A��L>�b���1��O�@���D!�*�������J.sQj7c��˜��ͷ^�Q��Y�3ٸ�0�"f����J탰z�h�g��&��k��Б-9%-���du�ty��	����y����/� �zG�p4f�z2�V�ㄗ>4L�KP0����@+?C�C#K6�=����sLs �nӳ1��'Q������Nq��
@ø�(b���Xb��gz<�˸�� M���a�2Qm�<���*ȚvK�<u�31�9�z��b��MP�b5��Mk��	*Isǋ
��_Cq��S��S�����da�~s{1�HǾ�8���*P؈��w�H��L�n�U|
�h\�?��� [G�G���T��p
W�!]��q����Ɏh�w��c�?d��t1��_���#������1�*���M.��׀q����0]8?j�Im)Zd��lT��r xKc0�䄂�A�g���{�%�}d\�;�b��q�sv�,�L@�9����薕�k�]�SrJ`�~�ԞV�HEo����4j�a3��AY��\k��Y>�Z�3�{�YG�o�|j��$���]��L�����������\s/b!&N�
~F`z��Aq��ܕ/�iꥉ��$N�7+\��,�$��V2u$�4*x��5z�y*��Y��� ���a������%�4�M��ew'�o��DTGx? �$V���YfB[#i^��.3�hs̟�l��.�>`%O�Z�V�_o�Ek�njچ\��P�xǔ�m�n����ޟ2��ț�O�8�,z�V�/��A\Km�p�I��Z.ov;����{�鰰�ǉl���S8�m�2��_�#r0O��U�e�`o�r�ԁ�4�xqC3����4�Q�S>�Ƶ�*�N�	y��-��h�K�g�֚��x���6��U� s��.w�?���54U/��9�i�SH��uD��סr��XOV��mT������CY�E���q/(��0XG/Q��e�g�/I#!�Wq癇Ӏ��6s0EQ�d/ՙd�"�7(�����.�+ٞ�l��I�1�J���B�f|�k��N`E�x�[��t#�kq_�9'��e#v���@6�����w=3J
�ZR\`ӸCS��I����H�h�~��#�
@��1��;U����5wW��D�pH���*�=����`T5Z�/�E�G�V�̹��4wVd�F�xg=�3��F��'�i7l,�|������h�,u1[�K���I����2���,?r4�l����KksW$�)M�O�*��(J�����BKЦ&�0��&�r�nˋw���O&����nZեV����G��
���חp���|��7'vA�\^�7�OKi���eKݧ�ȣ�C�<3s��yL$���2�}���+ ^�W��rK�
���s��y��6%Y�3����[ѯa�{G�%�Εs��+}?d�>+K.D�Ʈ6�h�Y��l�p��t��ӧ�����Y��]�h��ۆ�:a��4U�0'z�`Ʌ_HJL^�ā'�Q+�D��E�!jI�i{���mɻFk�=���8��b!��E7���f�g�ۨ�1��9{�WZ�[��'�B��;��]���,�}�w�f�2:�='�X׷׎!����M�Z���=�m�-��M�%�i���:M�`o���}1���zx5H����bޘ냖-(P����E5�)-I�G\�kE�+�m�M����#7���o/�J�=���P��N���x����sM/�,��z��9K���V
�iM��b�yz��Ƈ5����F��0?����e��i�ӫ�x�HC�d�H���%U <1��c�����V0�D���I�ʂ!�@�H�"�H�Ơ��������#K���Ψ�Xe���=jj�SXs�E����\"���̀ɥ��/fl؇d�(�B�@�1�p��m���U8-"*��~W~,5���N�J
��� ���m��-�5���P*z\͚���k�:��Z�rn�87W�^�ǧT�YQ0rn9����Ⱕ�"T��mh#?K��ZrJ��C\�S]���J���8���J>lI����Bۡ��)n6`B��iT.�Լ�v�g:��	9���D2�<I�fy�:	�f��0>�o!o�������p/��.����U����Ñv�����Œ�������SI�fV�����=ɷ~=rˤ���e�(��G&��0��r��4�p���T����4�'���rC��s})]GB�1i,n?߀��o�	�Ъo��{�vt��mcl��X�����r�D�y��돩߲"�~U�#Sߧ��c�Ϳ�}-l���u���n���)�Feq���t%�U���t�w"Y>�L�p�Q�(������Ai_��.HE-��_��[d�afCH�%d�,L^�uS�#L� �MD�������X��zt.�&X�*����i�Mj�f��r�aC6�%xk>�,�E�!��O ���w�O�S��t�U�� {��W����H病�é�ı�#�K�Y�i����A�*:&w���g�M�fom�'�C�S�I�s�G��DN�j=J�n���ޓ���x2��B̲�|E�H�FD�@�!���D[��6�o�#�!��ne�W����Ie�^j�Z���R��Bч,�4���}��S1G�C�G�%~/Wao`(z������g�ϴ�x%�����u,����� ~4�l��(��e3�E�6���Y�����~�H�n�P��b�:�!�u7m]ڋ&�U�ڙC��`� �x8��]v�}�� �/�>�K��ro����C8!z�j�5J	���0~^��Y�e�,���&�B&�9g����e`�3���M��,@ڰ�t�C`��Q����nb&kX[冣kv$!�X�����˽V�>�����'�m _�ûQ
p�*B
,�M����p�s��de������8i�����M�]��[]nC���и?7�m��K#"x�5u�0%2D�B��vy(���� �{�hw]����){(�"��w�D���K�����?Q�-�I��zܱ�WܤŦ#��"̏����GmKx��?�,�:+e�eKC��-�O#r���>�����S!��K�j@�N.S�$)F,�XQ����Tզ��u�Ƅ���?��n��v��uL
������JʝV4�J��.3�ݍ�۪-�����r�]�T[��z}Muc ́Bx���ˋ��k�p=��F��%H�j�'�?q�8'"Y���OZ��?ۥ0B��Gk<N��`�ʅ���-x�͗yL�FY/r�l��D��ӀC^��>��:�ܴ,u�#�)��n����������~��j`	QT��>te(�Hy��&�b����U���;��c���u����:7;�dU�X����L�@$�Ҟ����U��� �����KL%t��};�Ӡ�n�l^�x�&�j1UpÞv�RNAao���uS���5�jz��p�亂 �⸆A�Uހ�?�b���@��U�6L;D��/��5�Z��-+%�i�'�)c|y������(�g�$uEQk#�*\w`�9Ï������v;H�9p�Sd��h���d����[[��$z�9��`���2o�[ҙ/79�+F!h����t��(��x���且
>*F��[^ͳ�3:SHڴ���!�7����� �S羫�8�, ���
�KՓ�"K�XNsZ2P/1���,o���� n@�4^�����_`}3F׭�>Ũ�i�=|k����χ��d#�?�Z���n�L"[T��T#��2��,P����i��'kx ��`i
Jj�������&�����V-������W�2���r�Y�pa�>v���ǀ	�D�f��0����c����WO��I&]5���Τ*o&�X�qCC�m���\(X�"^ �?Uz�8K�+[��+b�Qg�`ϧ��&94&�P��VKd�i�Az�湮�(�5۲�
��"}�BYۺ�3�ȋ�:w�G9�*S��5�ARA�j'��B,������f�o��S@����~��#�FMު��+ǰ�C�D��PB�x�n��{������*,�Оs��Xo�Rx���_���Jr�ŭe�,�+�Mc�϶*�9�%�T�DѸoc@v`�!B�IH2�~2*�Zǽ���-��[to7@�K�����n�j՝�b4cWx�J�"�(%�����:�;��R�YϺj��6.cz�H@�� �kƪ�R8il�氮j5����,�T/�K��]��=T�M�	�d�%_;���5���:�G����'���M�*6���P�!����J�M�%Ji�HS��2g>�C������#�dD�q]5B��T�'w����e˷�;lgЭp�r��J�($}���,�K�Խ�Tũ����ok�.t�k�߉_����W�#��7 6+9:�UUdЊ�H��`���"&6D=�t�헄����1���)4��#�/�$�aW>���m��Z��K���O��|P��P"5�$?��Jr��/:��G��)	&P���W��X@���A�|_EO<O����z=�)��H�cE��A8��F�5'L?R	�+>`�s�ۼ�{4��H]�4pȥ�O���ө��m�������� ~��Z0���F+�I�l b%��C!�p�߷ׁwz w�E�c�ΉɌ{����ߴH�0i���B�K7N��p� �d�d�%���/B��C�J��s6����LrrUl��ǏVeE8U����dޒ*S�8�aܩ��\G 8/<�8����:�Þ���7���*�p�ʰ0+�I��
L�������K̴�~�b����؝�9�N���1�g�)	���s��9y~)�Ĺ�$�$&�Z��A^��n� ��8���_�K���Mgc������}2����C�e0u#B�*�0�dg�>�U��9T�5?"�\cΝ��,O�Q���������I�,]�O�A�	��c��	��ӳr�L#w��w�Z{��;�������yXd<�_5i�j`3l�Έ���F���k,�<��p�Aa\aς_���'��� Js
k�֮�o��j��}���E����K��7��V�� +SUbO��<zǑ���FJCu�MڜR��|���'�%	���&�@�������S��K���+*Fڊnw	.��K��H��-t8�״Μ�f\��<�q�����ʦqx�s@���E�w<;��|�����#��[o�_uK\Z���fδc	F�Si�Z��J6�����Tm���:$� .�'�c�@㚘i�mD^�@�q��g����`�!&!���N]|>�%�s�2~�� & �if�<!��C�>R�"���4K�f��[�*u��������>�Tu{��y 	���XP��c�)�����=���I����he]��f�c�����)0X�kp�L���l1>ĝ�lX�_�|����/��> ��\$��9��L�Z��y%��r@ �1S�^m���;㡠��s��/n���9� `����U󥷆�˯��Ӿ��.�@���<8��z�L$F>d�n-�!�$E_�]���Q�0,� ����^����fM���	�p�n��f���J���f\�!��uT�,�x�n�)�|K�n�9�K7��ia+�����o,��o��5O߽�(�9}�s�{�.vE8 Q�m$��K�̞ar{z��薿G����u%��+t�1����R��O��[�=�6<X����)��0���Ğs�j��������2 �)���Z}��&l��6;9J�����`E	n���7� �i�CFӣ�|y��G�3'y;��!����8�Ś1�s@�2WV�[� EU���
�n�v-/�2 ^��V��+�M�H��]jҠ4=؏�xŔR�)��������X�u��0u|�ſ<�n4���|a�=�^�Ӓ�)���6p!�jb�k{a�$,-*���1���C�߆]��>1K|�E"��QHM��n���`��b�>��t�b�i�_p��7*���n��w�t˞��aY�U����r��_[��!F�S܊�����8+��r�R�H�~�����Ĥ�/뮓"V�!cU���s��V�Z�]3#Y�s�B*I~�d�uHn�4�d-��NGd�1?o����n��Չ�d%�#�j�������i���iz�-�b���U���b�8�>�;jO�|U�����g�W���/ȎC��/XVٰ�]���ڵB�yz����`�~n?�z?Үm���~���y�5���`��భ�W�Gv$aɫ�j2�:8�	�^��˕a#�AQF>�=]e��y�r���Z��i��j���
6
�U�g)( @�z8u��3b	G;��8���I;6J�F�$�?*��ӈܸJ{���z�ɹ�D�C�K�/��k04��E����؃��]eNY���O�5xh��I����}'�@��%���l�n�\>`a'-�u��N�{�1���r}X��XR&��4:�h_�%[W�]��3�+Y����QA�*��Lz���O��^<?�˘�����(&�6��?+?�(sLgǽ�-���$�+�1�7쉮V�ʄ2B�]Ň�A�;��?�kP0�7�1���q`���T�b���N��m�Z�q�]r�nܻ�8��4Z=�y�$nu l}��䖪N}�vh�M���s:(�����'{���Ol)Ҩ����s�(CO���a�/�N�)t�4Py�7�i
r%���L�n�f���W��=^>��WV�X�w:�$W8��=mڏ��^Z)�P�50�m�����9d��@��հ�3�N�L/���ԡբw���Ӌ����be�J��r�׻)9��sT�c��L�j�Q�2�hn�h$T�#6=�>ޑ��s�g��k>�:�?�j�/	��6@J�`p����S�p���=��o��`�=���%�5�O��&���7�NUJ.�����he�?��49�U0s.<BgȦE-+W��#L�z�y1���1�FӾ�Ī�,��R�[����;�ICX��kxl�J�'j�7��H������J�O,������"E����P�%�%B��jv;�'E��]7��K���#9�_⥝�`�vk(�a�4����v">�X���JӚ�Rb@�����}k��W_��?M��{7'P�{8��d��`�>���o�1����"�Ω�G3�B�E���=�*�����iV����*Z�g����m��qZG�yȑ������+M����c$��&o�6�X�(�G���"Xp�'���8�oO��5�%�E �%wu�:x�y�L$I��᮰-����U�ӷF:���P~�}�`�sfih�Si�U-n�84���O΄szLI���:}�p�Q<Nx.�	���'�vԞ�v���V��!�װס��	Bd��}�cIA�|��H7�Ĺ��![�)��,'q�M�lֆ�����y^�@��prl��Q��fM�z)��xp��3H��ߧ#}��.�?�V��AQ�:XG؞�׀��W��>�U��[��'�1�]!�`JO��C��kv��Y�74i�,�GB)��KZ�$�Y�K~��ܭ]_� �ZM+�Ӗ�Z���]��L4a�g���C�î��j�(��������9+#~6�ug��g~Ě��5��a���:s����)�ho�+;K{J�W�A�Iq;{ �s�^"��ʰΨ��O�.���3Hs5቏���8m�lٓR?���8��  �`q�nd�A��q,�)�#�z�8:��oщ,v��ShT�ɍs����G$���U��un&��db-��-�9!�)��.�H!�~E��a�Ȇ����y�BQ06~i��^�E���ǛW4}��J��)��;��=�P�v��W�T�,�_O�mM��W�'���2��/�ސ=�j�tM�8���VK�;�/ҞQ�n���C�`�y�4�v���y@~cs5?����h���m\�!�n=��:�8���<u%�X���`��}l��.ԫ}x����:@7o�WBQ�k�U��,G�({�5�5�x�[V���ʲT3���
n� �z$!=
�Kս1�(i�5�{��U�ۺp�1�'�N
T�DZ��~�h[��kд�1��t�3�=5s%�LCU.2����
�w,���up��V�&l�������sI䏏�ܮ�_ύ�k��{[W3q��XlvH�6sm����_h���g�i��o�~��v���L�N��Si%��.��gѹ��x��zHOA�9�����a��[��Q�f%R��ksD���,R���);�cr8�{Z�f��D�B�w��.�+L��ǖ��Zd�K��l�:�Az���\z�ߜ:����p1z*��ԩ'���+��A��*����ռ9~@RZA�u�� �p`���$'��]�ߦ5�ĵJ�@KB�X<���/u.��Ci�:�G��+��P� ��Y&Z�A�ς�����⻶�*����d�d�	��*0��jyr�~P�t�*DƚkA�c���i��f�}�I�'0�ڤ��|�x�ϛV8��,���;|�]M�h͡y		��o�ԅ�զ�����n�Ѣw-����P2(i�|��������#.��Z�8�;�bpth��m�udF�I9�A�4
P��� �%J�g��u�������f9�ӹ���Q0l?Ae�ޔC��Y�P����i�����d��=e-�+�砍~C�.3�k{Eu��7��A�II��y�q�Z�1cڡ�o��#l�m�avz��,9U���PR�'��5����5PY2��v�����t(����u_��M�?��F*)Z��g =���G�Ut�c0���>f}��$�&�T�S,��t)��y%�}žh��1�Ls�x_<m��z����!O*�#s��2=�qr�}�'��b�<�f��F��N[1��{���H3x�����k�~����y`�9�utXvش��7��Y�O��VK�HF:\��tg�G�	�Mjes�q_V����W@�iV&v>�� |��f�g|��8e<�Wq�`�h������~t�nc�#Ť���rj����En�<k�x�<��������3�����9>5g���)$�]�H�١Z�9J͏e�'j!+��z�˨�"�SU��ٞ���}��v��v(��ر��P�I�Nv��hG�D���m}�G���{r�0�� sB�kSN�4t��G����y�b��ަ�"i�0	CČ��\8E�6�A�ħh��|�Jw2f �ܽK5vB�]��3'�������O����Uj,�M��ǊJ؀�/y~���X�&��?Ӷ֮M#����<�z���2�G`[�tܴ�������
|�����i�H���:U}�����Y��U�Bi�X���9�O�֯ʜ�O�Y�����4-#�`���e��3�h��5}{�H#M����� ��&��\:�����RK�f� m���WM����Xnތ׹:w><�i0��� �	п�yK�nga���y��&��r���W�4��&�-�(铯b�W�wag_f¾=��u�I}����� �����z��ϳJ��3�={���Cho�J8� h���ҬI����#��Uq6��R	2��)h��ߡ�|��qn����T�<���(���������A��9hɇ�ͻ�jUc���eG}�-m�����z���E�Ԇ}/~�$0r��҉8�z�&�����hB����?Qȶ^"���[����}v|U	W� �56�S�&�w��O��w�7sXi
[���{2#m9�1�������ǄJ�($�i~�����đ���?E��w$�%�c�q'Y�S��W�`0/(��1�"fD�a�1�6�t�=�@�,g����%�,�9T��6�Z'�Z�XS �b_�?���GbC��yx�je��J씋��T��X�X##LnY��~�Lft�����@���(�h&TϾ�$��Q�{������i��	�9��F�R��V��BLm-�,�%�ũL����="u�Ű7�� �	6m5��GQG�m[H�!�z��%収%N ���sA�D��/�-A�.�ﯟ�Ĥ��vs��k겹j܌ʉ_�����^+�dOKD�r(�[�ge�!eqN6�f9.'
D�I��Y�%�4�"�cE�v��{]I�4���7���o��~�"��|R�a���Q��$'�0�:�X��>o��p���P>(�d�5�8���@�O�>Z��'|����e:�<r�;q}��zA�Ӂ�Un�$�d{�VP �_�0��_�*��|�/~��<�q�dx��HW��`��Ŧ��{q�=��;��?��,�lm:q�}�Tif�f�ߴ�|o��\���ԪU���5E�Z�Ew����D E~��n���,:��GK/Q�����`�bfF�`����P�C9Jo����-5�v��ހZ�$������#vp����G��ڄ�Hce�CϿ���O-Iv�I�< �x�
1U�ګV�`{��v �J)_���\� 	 ă�f�O�M/\��#�)x�q� ��e���zN�m�P������xQp����\:�]�d�j�7��;�>�<し���7\��N�v.0�'_�#��H�#�J��rF���%�.���cj��
}�~C/?�V��i����<+�v�4W��h��b�h��&�IYn������:���Ԋ���,	�,��b~�Tcs���q�4����I� W��$��cg
�M�i޻��JW��;���h��x������2J�E�"rc��*�&�����/�
:�>���һ҅;L�ٙ̾�U�5ė�O��5��m&� M[�,v��WXX�J�*�(+hAQ^j�
�;�=�~p�����%�%`�{����Xu��%��PcwGhI�o��;�~]��ZĀ���CƱ*�VoVz��=B_ڐ�?I��S1T�f}2�%��7�G~Xc!�w�̖�/`l���I��O�����hl$����X����ǥG�]�,�}R�9;6���./�ѱ���F�M�
�\A�l4|�m����hQ�4�(�f��=/05{Z�{N7�K�ݍ���d�?�����	�����LR��2��b<�AcW�PF^�#$��E�x7s�T>�%�b6>:Fr������<�]�.[�5���>뻲�d�{�2�V�J�'*���ث_W��_������D��'��Es0�[(�����mQ� j�!v�1qߵ�s�*l�̕���[��OB$䍧��w�y�n�@��h�Y���,��wY�ƾw�s�2��24vҤ�~ة��.�r�_�6��S.mX߉���5_vLQk����#�'L�(k�_{��(P�9hd�Z�՜�P��R��	e��0��n�������[����$�9�"�8�Q�X���֚+��&��J{4$�7^��+��&�K�=��_l���E����{c���uz⻜ڞP�{��IB��������k6;<&��e@��s�̤Mq8p��Rը�/6�I���ߩco|��5�qՌ����a\w6;�� ���ul�m �������p�i�	@4�U��0��w7������H�ۯ����Vs����e�B�Cg�=��-b�\O;~�jN7G��$_��c�)0Uy}���-R^�%꾮A�������D/�R�6� S�e�:vj9*�yc�c��`%n��K�(Kz�nb�ȡ�9C�� �Ϸ��x��:}g�{�
���/O�ǜ���b3˅qo�[�P"�dr����֗��sZ�������#'��R��Y�~����l�e.D���.4���K-�zėc�>�ulX4��@d9u)�\Ph�{h���#�#��r(QI�ꈰ�D��a=[s����7�#����v�6=A�d�!d��I���WW΅��	@����D�|�� n����[������Y���/��W+���{k��=A�RGdAܖ+�~h�OPZ����@�W#+"6�qig�b쇘�-���:'�>�>OL녷f�(�-�s��=���<B
�*��5�8>JX�C@�Q�x�kt�%�8e�0`�3-)�_���ûπ}�);��h��w�Y�iu۾����/g��R^~>��(T�iۗ�Δ��υg�a��q�������O��y�SO�۱�|����}@��~�IrO��2����xA~���}�U2s� ��������x��Mp��b+���փq��t.�YZ@����x�"���d� hR)<�ߋ�.^�N, e���e�x�;˭��O���Fv�4
����q�u�S�>t=�Z~0�����>��O������	s����J0m~Z�eK�R{�xkƂ#5b�<�UК����gޒ���|�}�w������OF����v�9�e�=���93����!�xn,c"���C������H_E� y_����7w
�g�80��!̓��F�^�54���8�����.*���!��{�������Y��n�� R/�Y���M��ε���W���{k����4`-�Y
�;XZ<+��v��f׭�7!��Ad�T����r��D6��b���i�M�5�Odz�A.C _9�P�ν�Bp�q`
.�R�n�p�L5���vJ�Ez3���9��oeEe1���>&/�qJ\~����m���jdb������_�[ʴpQ��1R���M��Ϙ~��:�q�����3^�A{A8��G%H?,�O;z誱��в��hf��sm�u�����v��2~@]�,��_��a#Zǚ�)o�q��Y;�a��h��
���qVK+Yz��u�c�쫡P;~�=�`!$�]�T�#�0����QV�Ȓ��2�o4f�p
O�'�]�`�C$�����,Q`�0�g���:>���K��pj�o׫��g� x$�_/��XB<�;�zjP��&�(,ë/V�p���f��)¸�H[��(�]E����N|�jck�~")Z���-:MiD�[���7�h���Nx��A����m$��U�{���Kȋ�+G�^!�-��^-��c�7�
��cQڼ9�v�>�W:�o�w���P�J#�6BQ�I0���@DN6ʱyr�;�}�~���n+�`Of��
'=KE_a?���,��̤��]����!97%?"�H1_�w<�7�Tck1ehMu�g��f�?���ׁ`�Bf�i�zFigu7>$�T�Y'���&�7J$�U�K`єO����!�/;h�k�k2hp��Vd�$�-�{�qΰ
lw%�hrܙ��?ϟx�:�����T?�Dw�J�I$qyim��SR?��������JV2�Rf5B��^vԤ�d���)"�{�,�R�
�Ĕ�a�(����?W}��l���-��׼��D9��r�`T�68���8nPvǭ��Ն�[e����#Y��.���@�NX����_�]���������w4���k!}	��-̢��i"q$,��
�ks�C�HJ;���(j������a�l �� �X��@�/-o�` �>}����!���K���CW�_ռ�= ��_�q����[��p�<����q*��*+;���G�L�H�`NJhh{�4�D��`��.�n�ᑭy�ʃ��E?a�?o�JD��,��8�C���.Q�2q����#L������9�\:�� � ���JJP���,	�ml-�u�ܲ���0��|��dE]�ݱ�S>gk�S�e�r�!B��K���Y�z���T=^�d�̀��ޘ�<��{8"�S�qgs���U����&G����Lg�
���,�mP��7:��ćԣ��y��fS��w�珫4�=�g?��{c\����P���������������F�	�6�E���/���'\��$y�<"����b�}� z�*��Qw%("���FB2Ѷ]'�rm�8c���������g�v<�_vm���_���;�~��2hG�wW�;:���VeΕ�.*�t.����E$GH��_�h�UU���pWn���q>�<��9���������h��-=-��p�PHR�iJL�X3�)l�5l��Ci�}ڞg��i ��h��!�}���ml�����'��ȓ�%��yS������n$�H����lB"j�w�5z<p���y#Q�s+ӟ����עX۟%|�D��Q�e�ZS�'lSͫ_a�0�N��몼_��,[ <b�oE�T�{�x�����$��ݮy^j�C���,�Q;c�E�ǻ|h�u��K��6*0�N
|ϧbg8#_b���_��1��K�*2�eE��PY�F'���?Ɵߌ��;�7Vݜo	=��%�����Ɉ_�F�?�K����PN[�/��yY߮i>1&�����ȍ�D<��{��n���)�S]�7�`o�Y�ē����G[�E5,���oTA�����'�174>���8
|���Z��D3�w�Z �x�S���."H�?�S��|����(�� ?�e��3�E}J����k�s�+�!�A�$\�Ļ:n����_�O'3��LR�0����q��Ɉ������5Ζ@������OW��'�D�Ƶ�g�	ޣ
+\M�c����ꏪ�ܼ �m�i0	�qm ���p(jv�J�n4���>�_�D��<����ڦ~TL3�[Zф=v� ͧ��1�s���M��"h�[��iCv�2� ��̐[(j|�v��f�������[�O��O��?oX�z3K�q���U�����+��e0��N�Ů��g���0�
~ָ]=���̈́��X�B(x�!��5"�bK�<����:+�l/�x)i�����a��|�q��[������wt�Wn��l�,R������7ߡ,_-چ�Ǉ"�3<�8I��q/;A��9E#6G	��?��C�൨\��I�	�=B��C��h<b�p.� �������}�~O�D���~4Y�gU�t��̼�%0/�}¥�j/�3�aڋ�Ɵ�Fh;��p3�}�9�$�qo�3Ee����I��nlp�:�K�%.�I����F��R��K�} ޣ9��a�6�B���CQ�/8`d�V�m��C�/�dEd;����+~�K!�\���M��wu���߫v8g��~O`�>å���8�����RZ�]=��s�$\�)��"h�ۊ�"p���J]��V��?b�����öH�wj����|ޝ6M�yנ�nq�OoB�'tƾO;��X��^^�@O&yh��껦�}�����Ls��2�>�~�!g���H�Z?��#f�t������rX�����wst+*H��]��./I?��b!�=�i�{z�7?��2x�<��سz�y����l .�������:�Wݮ�;}�Q��Do(�u���tU�~z?/�p.pz2�9)�oT���MR�|5�'+��,b#�J�}_���`ܶ:s��!p��*�xȀ�к�O�M��\C�uk�lξ�>��>���-D��F��M��\L,h��%Ǳ/W��z��GE�m������=�@�/�(l0>l����
��-��.��B=���v�
��\���qA��v�u�\f�o�s$R�<PO�QEĵx^�Ba ��7����t�����IN����n�m/��Y�K�0�s�*��?ɸ��+��=��Z��|�m]k3�
���L�#|�o�;IT��)���	PDţH4[�����!ۃ�-l��W\*)�����EsQ �Q�gT��flG�:K��5�ٰ�����f�W
��99ݡ�㳂���;��5q6lo4<h��X�xy�|���IWttU��g:�6X!�!�|��V�oz��񃃭쐷̹StA�An�9!r%\�0����X�����7�?�.YAC������${�Y����֗�]�<k�/{� "ȇ]��������rf��n\�>dnK< V�79��|e��x��kf+\���^���������8	L��.N����@�Ά��j�jԼj�|�g�8C�d��k�\���u�U�fi�$��˂��mJM�������B�*�_�I�k�i`��@	wIx�&W��
.m���2��Y!���u"��p���Uy�QH��S�p@_�b8��ò����Ơ���a���pCP`9w�xµ�2xq0�PAP�P�rL3��X�{��>a�A��yF����B @����0���NAX���f����X@ğ��~���)҉b�*�xA�������@�(�|nɹ�wE��+���e�S���&��{��,8zeo�Y�1Y'C�iv�:~�l>5��E£���7��/�^�?��r��\j� ����nuU��CN&����M83�����t�����,JݧU�(Hg�aL�� ��3ր���,+�GE��8�	g��蘻���~^���\4��V�B�Vs3h�ؒ�{4D]�����~�u�5�?B7�e���Q�&�V$%¤��^{�n��#8�5��w�{TYG�5@T�\��x3�&���@o�vӕɽ�C�X\�����I��2p3�g�v������z�C�Gx��������x(S�4���I�2�tU�����C\��8P����U��k��6e%cTSߊ�@�:^�V0?yQ�3d�j���*V�v�Wbǒ#N�J�Ëf��z��h�(���"� z�]��C��x��C�3C�
%��XH����R~��B�r��#�_kHi���͂���N�I�W�c�ö��c����t����~�T
�Io:s7�_8>z�[,�'���0������ѵ��A����C ��ZQ�jc��(��8�;y2//S+CL�W�"�hYu϶����<b�)���!�92(�&����A	ꍐ����w����?;,���w�J0����8���pw�/�R��В9��`��k	X�W�� ��X+%^s��J��^�u�c�=��p���rL�ڻ�	�x$�V#S�f��Nso0��I�]%^�/��V_~��ƜYA��c�Wz��WFf<���E¨�z�+D)��Ѷ�z�
���:$����K��`@	9���$��)��]�@��Q�]-&�
�6m�Y�"J)�\�V�;cP��j��t�����~��	ń��-SC��z'B��	=�.*���̋?d��Ѵ�=�x�?���ת #�*c��s��~�m8�R`fF��n�ڸ���L?�^Fh1�}~�nQ�+.�o�V��X;�
�~�{��4�.��P#PD	��������E��W��s!�3��Xj˫��O�^���VB(pOX�i f�Ogu���Q���3`޺�	�7$����)�e��L8�1D{:�=�!z���ۉpyx݂k9���a�V얿�:_y٣nY�&r3�A/��}L��b�l�5L���ܣ��FEJ()_�L���x!�^s��c�	�lM��Zg�� U<�y����P%��F�l�s�+\,�+1�AX!c��*�V5H�I��UG0T1-`L<���?��̜��ʇ�ŕ��JUXv�I`���~AX�%���&��i���_��za�MP-���)0�S�t�0-2����(Ͻ̅�}��J6�#�5x�/�)tL�������ߣ���]�,��_x�qW��b4�&��t�C��{�#�ZP<�d��u��$���Ǥ��x�k����=���9e�i~1�uƄ)s���C�i��;���,�+�;�UO"M�ũ� }Q�o�p���FTB�I�җ���,$lf����z�d4އ� ��K���pB�n��]|���;#�Lܧ5��1T���E��t�d�]~i����Ɍ�]����� ;cЎ*)4�t���U��u�>�U'�T�#����G;#����{Cŝ؛���F��v����ڡ1�:������G��+�$�����dB�|�wU¸e��^j_��=ظj��^�" ��ƛ3�2�p%5����oc ڡ5�Q���uΌSͦ�'{u���rT�҉����u2yCY��o�i�W��>��8���l}����S,��{�GE�&]���X�6G���/Ҩ�*Y���'��jAk��M0��h0�����_+C��+j���V�P�����8���b'�I�D�~�����$������T�r�Ԫ2�V!��ΰ ݲ�`�����ŠO�4�]N�˸h\��"�L�^�n�U+v�r�����٭'#�M�QW[�����N%\ߒ�)�S��א5p���#��O�K�_q�}�W�"
���7X��=�S�p�4��%k&?�6Ƌ<@����n7��D������ɱwA�ь��Ļ����FɃ�����B�yPM+.����a�2R=�������3aJh�K8��+�3l�=a�k�r8��r"��J�4%>�#<�27Z�{7���(*z�F��w�K���0͐�񠙈'��$��%Ϻ{��1�t�`aĉM�UW9�7�"����r�ʰW��SF1�
��z�L7:�ק̩��p��\ί���n��~B?H_�>��A!��ר�b�+d�ʝ?�`u���K��I��\J;)����#���1�P�;�����J��	�xh�<���9F̓� �ƏC$���~`��(�Y�:���Gme�-��l�X>A�
���˖@FrbQTj/�U�z�k��{��^�C��C~1$�&L��Jܠ!8�����:�� ˴�)6;۬6F�>���*3m7c5�J�«�M����D��� �ǠMh}�-P��5H�����\�C�R�b�Dh��Gt��h��YϺ׍��WV����^8�Wӌ��{`a�Y�<�'f�!s$=Ȳ��ކ�N:��\r׃HA�,���+8��eF�?��T#���� ��y��Q�C{I�qM~Y������;�~'*���*Ƨ��#�J��f�"�\��7s�<�b�����*Ċ���}}�}��-R����&�)�L�)4o�By�dUI)xB�����,zĔ�*p�C �8�1��>�]��Y�Խ��i��MJ5z�����
L�_,�n�wPj"r̤�����&�83�c��݆�Y� ��t�i�3����,�veu��
8(�0"�!Kx!���2����/��p:�3��n0��=¯	��X3�w��*_m6������bo��n4�.$o:뇶eQ+�V�N\�-gHջS��
d���s�*��V�pa*qv�T��j��%��n��m;��H���J����c	�T2#Fb�,g�/�Kڡu�g i��v_�Md/ac�q���r�uED��>W$R�hı)�}b����3f�am�h#6T�دt�p���I����z����������lg�l�874G_�3����}N矮.Y����9�n�-�m����kjB2�lûsj?n�����+�Su���N2�zS������`���v��S�v��*�
�M��	|���j5�K���{0��� -5���]�<�beo5)�^j99:O�ژC�0��P��x#P��SiC>w;�D͎׉��+R��}�x栦����`�<mlZBZ�h��"��i r	�t�������QC�$�|��.6h�O�Y�rZt���XJ�n7�"�%��pO� �����������OG��R֖���Z��(o3��}8&\H(�A���c��p���]�ȇ�xޤ����7<)�B�f>�������pNXY>���f�P*�ct���E��q�2�%��#_T�́e�2��+
IwCoˊ9EJY�D�C��m��x�o�n�R��S�kb.�X[E�}�(o�h�a�i#����=4�o�r��_z�����4ܡY�n����i}��-�䕯��iv��؀B�5C�\�B����W�e<	ot���� �w��7��c�p��C�d��b�b~�V{�BH*Fr�+p��a&�b�׼�D�C��=�m\Sc��Y`��Jt�Ȩ;�إ~4�d�9.�`��%���\�� U����o���I�#t��Аǜ�4��3��I�"|��+�����D^��O&�A�&M�}e>(Qdd��ŕ�����V���I��^� ��@F�ʈ�PY��c�����:u�ZT*m+>m�PO(�e'�,Z@�4/���k2�at#����4��b���s .�n����e��DV��рV��1S
T3X�1rn����	
8G݇�K��ݜ\j�~u�Gog �~;R�Ud���b���2�8�
�|�Jѭ�T�����맧E���̔��w��@
&0N+JI��L�I�$�������ɑVp�uc��#�P���2�E����%;P9{�إ1wKo�����#lĘ�:�J$�z4i^si>�J�$�N����F[B��T#Dm����;�R�|��:��=���ù��d�y�]�N}��t8˔D6+^<B�6Q��nM���uVf</�� f������(��~�Y��!E�oK_�|����D?�p�!6~�^H�f����۵���쯖��;c�(���ћ4�l(��O,�'O��5����s~�+�j�"X���F��bgr��+Ϻl���c�f���`�8׎{ӏ������N��o�����_�sU�7��k�p'ۥs,hz�N��sY�hRr*����"+���P,x1�m�����>���,`N_~�ix`H|��� E!.ײ��V����P���/*B��
eO�����w����{����([K����v�S	V��X��+���FS��og/%��Uj��(�:��;�O�V�~�[�-@��gUe�#�M����[�SF�t�)kA�J����vjE�@��N�iEE�p� gd�0�H{��a�j=�+�v'��ky
V^�C�{�3��a���X�^,ךi!݉ݭ��&�Z�V���w��Z��{j�k�������e�4b��+�vt�Vc��wZ���nwwf������Ƭ�U��ꇯ�k�c~��>d���+���{q:�)u5�{T3�m�(�)nK�hz� ���� ���U�G�S�/ZP:�䔨o/SE���
����Rh��,z!7��R W��D�������Pi.8h�����Ѧ�h��T(����Г|ʋ��Ϗ��l�P���n~_]_U�}�XL_���a���3n�k�3.E��'�@ikwb���7��*2|���[pq&Y��P�/D���6H}b��A�`���/�ج:k��ORG�p{6�z�홨Y^8A���>%�"IO�����Q��o���x�Yr�M�) j�@2��6��cs���3t+a�u�u 9��e5xw%Eq,IDӻ�ʗ{4�����a�Y�����ߚ:���s�?柢�ED<T�+����Z��A����D���;
���^�J���B��~�{���R8LM΁I�f� Fݨ�d���IMЋ��Ӊ�=Eڶ7d��R�s1]8�U3��Cq�,��"/���Y3��W5le#��HK�@O����Z�:��/yt�/�o�6��4�KV�Q�&���*�|�kc1v�~�<T���]/�R�y�׼�uC��Ib�VH�埆�
��gPc`��ȘS�WM= �a�|���|4֪�F�٢,�|�"5��̑����_l"	���<Q
w��<}�Vf��*���:m���im����v��c�I��A����:{P6	�����o�B� ��&Vc�I�&�Rv/�@Gx?���̦@�9��ף�F��J�_�=�s�R E���Kv~t	�z��	����(�
��z���9��ZpY��ӿ�mK?��`M�E�z�� k�.�(D ���>���:�X��%�v���b��[.¤+�~&n�?��<���<�櫙��T�*��c�����c�Ei.��܏P���q���N�7r���o�{NQ	>����/{��>��5����mՐZ�	��SK��$�
T�	e�����4��H�U�"��H�lV�2oE[��Ka��c�*}pfCױ�Au�}�AZ�^#!���@��˴����-罍ܜ�z��l��^�2�b���E�����2y�n�� j�C�:�o��Zs�qvFۏ�vOe2�,V0P��F~z�f(
���Nl*��B�Dڳʬ��Y*0� �˼eĲ�Z��
��p о�=d("�-���@(���w�����G��AD�����z�)5,�"8�s6���R"sG�a뀱@�� 5�%i�����U��l���@���y�tN�v[���q����q,<@�gw��N�B���t��TMV�2�ڌLn�x�tݗ���1�Oytc��Z���,Xy���l��-��y~�K� �2eV���e�ۧ���<��OU���4����/�������Ս�� v��m�o��������0�����DT"Ջ���z�}RD�p�F,�qm�2A[�S,å����f�{9|��1��}��֕��ڦriv�������dQoנ��Md���x1HB�����@Ӆ�$ŧ�e��s��\��Y���C�����$X`>M^�Q�NՆ�c^�A;%u>�F�n�l�O;.'�� ��D��JtIA<��)τ�L�!~&Ew殍k�r�Όҽ�"��bG����+X�Iş.܀��:%�����4�<%��*�5������s��=`�y�Ob󚖄��.�t�c�)�����K2�F����<�$�[���N�%KO��g�.��\,��]�k�517�te���5��ח)M�@�Y���?�w�h��{mHIn����(��?C;?��ZC�Z9�9�I�K�C�``ǖ�M>7���	�[���=�rϮ�=���cB�V�oq-x[蘛���m��K�ܒ�^�f���0��~8��N�V�O��%Μ��{���0����q�X��vy�J��S���ٝ�I�5��ɝSoI��Z� �˫Pl�֮����6mā�u@�e�ش���E��

k�7����?���&�L���;�u|�"f�4��'7�1���Np���A�/���v*_��m9p[����)7����7�rǝ�K6���K����.���nD�O�!$��?e�J>�a���l2_͓�)�p�W���3�V�r���;^� a�����j�4"ݠ��z����z�;p�XLV�J]�����D���%��9�Q���^:�m��\[K��,3J�_�R �B��c5<Wm�z�����n��F��%��c��u�ڋ�r�f�"�U� �+�)Ȓct��2F�Y� բv@�v�SZ �;�	��&mC�v��/����b;�����0�����w^���x� tl�Ϣ��$�wc'��s�����q���Py����Ij�'�)՚�����w�u!�َD� j5��L�04��W� \�����ɣe����!ʃ���x�Pt;¢�~8(�Fa[X
ތ�-��0J4+��j�n@R��d��?��;�D��ݤ@9!�89N��Y8�����y�@ё���3�yHI�h%�-�@��1�Q�Ա��M���tFtݱ���]��-�)�^Z���{BE4�%V�9�F���L����f��0�i�7�rJ%ܳ��h�W���)�ؒm���M�P�6H�#([�7b�%+��++e���������1-��^����{2�i$�g[.�٥���ǚ�(�<f�[�c��!A��Xԁ�u�v&��r� ��\'����%+
<�|�D�l�����?�{�le/�����Dl��J�S�_iO)91��Me>�,�K�!
e]<ړy\�=��W4�6��my[utDQ��}6���Y���
�:,B�I7PS�r�l��CzS� �s��-�q��(^��s���8e;�Ȫ?0�%�juУ����*��<e�6l������3���Z�m�z�mN�s��C���W�p
����k�Ȼ�\���ܵ�&�����6�7"�fG��U�;�\՘U�"I�juo��yz�������.2�`vrJ�(���L�+�1<���1�UuQ�3��J+��b�.��z�����[��Dk���F���H���jN?#t/-b�}�Z�5� o���"&#%圂|��.rt�dޔ�)���r���9Ѓpq���k*���Xb��U{���lc=Tg"�wH�mp��tnP�T3|]ip�P��/�\(J�����	�.�h�m�U��hqM�O�%XJ��d�B����T_���?�������+y~��{��Q���,Ob"����Jc��R+x��rR0���'����`#֣�ېy�(Z7�����������?�Jo�TF�얁f�I=��߀�Og�V}?��-�U�%[����X��-������Dl0l!�6�=)��~,ѨEǊza�M���]�݈���c�J���0��~��VE�a�M���Y>k�������n��@���T�9>SR#�e'1��O^ND�Ҽ�L�]S�Q@F6�|�W�۷je|�E�YE^q� ���E���n$���χY��O�. tc�)�~����5�^���%��f4근@�i��U�v���khh� UG����|s4�3,m����i�����%h���nlb�
���|�F��j�krh^E
�F�ˇF�gg����X��� +Q���hh+LW����6c���7ܰ���b���zQ��KG��%��Mt�JP��/᫬}�"��؈Z�����c(�����q�D�ccy=[np#��C������������@��ӛ���)��&E��\���.�5�@��H���b
!9�=���E¦Z�a���� �!ǡ�8�(a>y�{>��|SD6�`kTd���\�5
5�-.x�F��˷���+U^���G��9���}4��gj
?'lV�`\@S鏈�g��ʞK^�Ń�(4�%����6X���.��韑��%m*>~h����9-":���fj#N&��@���T��qc���H��k����u��9��Vҹ����Fγ��`-�L�K�H� ��t�Jg��)��vNG�K����[�b�ͦ@l�Z��f�|��w�D��x�]X6�f�ި��ęk�ɗu��5�*�+�N x�����k��["�4U&������~���Ş?�5}�����.jV�`(凷��
���>�Q-R���Tie�KU���	�Lfk�)o*�S~0��W�4�Q�#����(�1��]��o�+
Tŉ�P�;��$����RjL0���x��ƌ ���+a���:
X@��5F�,�Je���͉�	�52�;PZ=9��M�nQ`w�_dU(
N٥48mhu���}�l�),h[�=�D����'�.�:O�[�_x�	Ѽ�Fd��>
V�hi$]h�
��IJ"�O�s�*e�lJU6]V�Iֆ{3�q��1�	�1?*N�M�-ȝfؑ�����,���{�X��INq`ɿKJcKXɲ�,U\r�K�������'P�_̴��9�ɑ2��]���s�y�V�;�:a�3�b_�҄��h�#�[���� 6\������QB_ҍ�Y<�ˑ� ��l;����8o�V�D9q�5[V(��q��>�t�V&��;0�I}y ��#��E޲����>���8l��N4���+��⼀�C'����e�E���"�����V��6�x��Mr�������a������w�M�h"S�n��C=ǡ븨�$��T*I �q���!{��O�@��A� ��߮k6�5׻������,W�9f"U��,35OL�H*�=K�DQ�r'��y�����+���N4��[��.$�-ᖪ���5������2�&xk�3s��_��
 0�����u��ɱ�^��VfgQ�
���Z���)V4�ԇ��6a�[x��������W1&�|t~{��=\ ��������g�7�jF�^�d��v=�zC��������7e�GI.�,%�q�T@E���q�j/>��i�4�|q�jN�j+�&�5�҃܌�vo.��H϶��k�۾���Ѵ�N�遏��-\ Ë�����j}Ȩ# p)G+�y�J�xMS 3��1�Z${׳z��FLx�8���i;')�24s���]sz�6��˫�L!�P�6(�$�w�s� �������zM���=�]f� �w[��XP0'.=эDno�d�PeapE�$����#��^H������N'	�'}���qƇ��렦���Z��en��S6?���=�'�P��.��v��鿴���p,���m���ɲ+O�u��B>E_�:J���@���p8�A��DW��+�)���0Y�R����jϯ��gO�!�	Mلm�h�p�m��9
w}nHϩbJIl���ǅt���Õ������#V�}���]/�t���]qX��S�yY��u���7�S4�;��X�ͱ�j�������� CC�Ǉ�{�?����X֦���k�T%�m�����[���"�x"�Ȧ�
�a����,�*��N��J��}`��LvEy��:����Ե���1.h��;�@��C�y(]#i�D����ig����-�[�o��a�%�~��Y�V@E��p�ǖl
7�:�x�=���`�2]�HY����4�S��}��t�Vs8�������������ƚ�3<���m��0D�6qi�X� ԪrVz�e�}t"N�а��	p�uf�A?\g��f,
 ƚ��M�f�i�1T�)��,�QZ�K���cԠ�c�2����}�k�s����S9�X�`���r[|K��O�_(�f���皆�$G���_lz:�L��>\)��)M�����U��m-N�+;�W��$(,?o�F�!Pw��lg�GXH�|8�����]�׼R�H���縣�n0���@���PU~5�R"�9��y9�ǃ9RdU���x�3+�4���Ú�xRK]�:O�����2�q����+:�������
I-܍n�}�Ϲn��ڿy6���z�n9!ؾ¢��)�Q�8f�ɹe	M�Y���d(�6����#3�.>D�QA^�z���>$R��R;�g=b���gS}523���q�fv��pt��O��X	��~nr�.�P"PN�5}���VmF�)v1l9DU(��F�/��P�������<`ر��}?����o}3��82�wn�b�/R����R2��Y�n�Y�� �k��d�qT�N	�/���僝a��!�9�+A� 0}�0[[Z,F��Y�l����*�����[��1|�U�?Ȣ���$^��ݨJF�A�̃q�݈�,N��Q�ʃ��k�9r����Ev\4� AR���'�n@~g����'NBj�i��f�&�(�u�dF�2`La��+CX	�	e�׮�'�W���N\�d��׼1��bχ�s�����6OEx���jްƟڨs�Q���aD{�}�x ��;��T��ȶ�X��v8~#��21	Rӽ5���!ҿ��QA�e&Q5�L���LTސ��l�}|9@Ɣ�e���T��!�'28!���&�{1x*}<��)Q|$�F�:�!\�}L��"��McDW�ia�\��C�[f֭�Ar�0�WN��G��~>���[W(�5�=ВJ�E�%����j�Ķ<���?��������p^�g���d��� �F#On�;��|5I^W���O8*p�JH	��O�Rf�I}xF)�JyԿǀ'c�̿^�g0iS	\Z#A�a2���s����;���%��q$�𝍢����yN���>?��n�q��y)��f�Q��'b��u���7�I������`M��+B�˔��
g?T��Ε�Z=�Y�mӅ�D�p~߇�k��yfW͹]WkA��iX*�sį�\�T�P�ڛ�&�s�7Yޱ w���SBN���}{=	��*�k�2`!���ƶP�NpNx�΂�;v�<m���K\�e����Ky+i����9�7!gf�Ƣ��p�����\�f�sW��V�6���oӪ��Y�_#W3��A�W�i�O7������5Xv �Q`Z,���~O� �����/G%�T�����$~��l��.�r���q�w�%u����-n���d>��vHǑC�y��zR��!��b�gfb�M�Z�{k�'���þL�*V�{囁#NQ�ɯUg��	8n�����U��x;�&����a�q�i�K��Ӓx�P�;D��}%6C���_Ϸ�\��r/K��uo�C�[�Ũ���'��9.��.m�''i�/b���c;��X6�#�8"ݘ� ��oՎ��\cD�J�CY�S����Rъ���ݛU[k�-�Rf��B^F�w��x|�I���v:�j�/}:����Yw*�5w��o\QC�\Cq>�?��Ui4�ϖs�.��6.j<Ȃe1���N��!Hφ�F̈�L۫���|��C��D�)ȓ*��5QB����+�+.UƜԠ"Q+�.��䋜	4Jd-��_�v�)X�Q�Z+�XfGr@�EO�&6����iJR��S��;C:�����H�t'�V ����s��apg�d���8m���*�m���t��'��G9����˪:�5	��t@VnB����y@���<�Nμ ���C��*�3O+i�����?�IקhQ����;���6��W�1����'!7���3J���^3ܿA�H��n*A�!>���ExE�QU��]�x�&�5��5�"�����O��� N:�Ik��jfk�Sj�E��&��ޕ��W����	7��@�4��`X�p�O�f�c�LȈ�s�AT�ě�㊽�F�ϖ[���sa���j���]���\��"�[���R���U�tv��>1��l�Ux�
�R���c�}k�d��;�1�]�<�S��f�:�w6�WQz	v/Z+�6=�,�ޫ|�f�⢦�)a+�o����p�k��2҅eH�f XP�Cg��U�Vк����&Q0
<ř�6[���7�e�&��Qץ��A��,����[>�;���+`�e��	A�iE�d�U�뱌^ƼI��V@Vd�8���=I�)I�px*r����qA�0Ͱw��?f�b�y8�Y�:cG1f�vȿs�	��Gj�n��w�'�H�C6�lݵ���v��7�W�]T�����`k�<����9�Y&r�V69�����ٚ�c���6a��U�?e7�1L�<4Z#	K�Y`�I�E�v$nL�h��jT��ϊ�Yd(Tӹ_�`y]�3��V�8�c�c���α���J�n�6�c�Taɦ]ѬҲIh��[Oz��*;�v���@��*U3�E�e����Q2^������*��ȱ%9�8�����?p�ۻ���M��	y��*j7t4�L|<��13����p�1f�z��z\{��_��9�W�!�������q�|C��j�k��u�Jj���3yֺ�k��'E^��)����8L@�ܱA��3+��弘ۥ<
D����~1r*b�}�c \P�Bb�ќ83��Οlq����x�N7Y�z�}R�s�,�F���V��R�6�D��-W5Q&n�f$<'�HH&t,_�W�A'�T�?^x�!�_���N�ݨeR8��r�X�]�$�H�#k�A�q��h=�O@�zS�_�T(�*�O�Q�-_�,!�L��Sh�T��R[��?,[ms�̹h}N�e���6�@��I�n� ܭ�4D��'��&��oV@#�v�s#���x��8)1����,��r�A
��a�_���2�m��f����g㯠�L=�7
¹�#aPCO�{�/�"nI]��]]�E�rT6��r4"P��f|��&o��k�?�T���h$_�PD�p���LnU�V[�����J�2�~�St�F���6j�zxwZ����do��;W(��Th��	z��"�^`����<�X�Z��f9"���v5\�?�E��6!h�-ŕ���G�qI�.tl ������v!K�e�h�NpD�h(�R�;�
h�QF���B��+�ք��FW�]x��È��Y��lkթ�ԥa��0�yz�a�j\�}L�v����u��
R���d��y�Iy�A�{� Y�mEp�Y:��,Ђg��m�
��p4�1�G� <_���⌍��zh���A���SnL)nUj:��tON�������>��B9-�~F��7�U�i���'�Q�!�G<�����y�������d�߰����PYG�\��漓),�+rJf��W�m�Y���)��q�o��l��;T�gR�����i�8�so�=���� �o�ѱV��\lm�N�h��A,�C��$�{�v�;�0�;�@iI�e��r�����h�w����s�,��̈e�����V�%$Sq�>{ob���  �;��8��K����Ōa�B��1î�A������>%�;dHD�j�����yo��l�q�_�Ļq� ^nA�?��4��Fq ��ּס�b	�8�.)	\�d���.���PP��zlQfC�-H	C�w��jMF�����/���t��nl���� Y�6��l�g�bi��h���^_�'/b*��<Rִ�P�=X�� nS=���(6K4`�v�i�w�#	����?��$�Z���N1�E��"�������3�l#s���X�OW�o^�z������ܽ*\J�oo;�7%��o��2S�䥛�*�����ˣ��ê1y�	�&C*���x�kk�1��]'sg$j"(���hq㍢J��[dk�3_�We��T���<	e�����͊���[#_��	�1�`�����p:M��=n�r��Ӕ��'!���v�8
�r$��-v�SVw�Gق\x�c���)��� �h8o{P��w����� ��+��]�_�N��>���(�fѾ�D�y��MU	����*c�|&�Ѹ��`���r�����<y��
��z�B��qp��/��ޞ�������-O���+�9M�*d-�������
r2�/���[]d?�+m�L�Л�A֗Z���f뤡 Z ���}�;C��뷟��J��r�� ��]��oc7�n���`}��%�����R�K&�����鲀��㾽yBaOQ��͐� ��%"2%����Lr�Vi���!���nu�i$3"�ڰ[p"έu.���X�H����$s(%il��GR���@i'���9	��� ���z��:���h)��^�
���O���qvT���Z�˷�Ym�4 79z�`nj�w�M>%����E|��R�׾Q��ni%
�/��e���Z(��]�J%��F� ��W�Y'��B]�B�MǩHLQ�� DI�'82d�|uy�b��U6��I�sp��p��K�gkŞ�w�F���R��ߥ�@Y�:Tb3�"�������sW�,�ʓ~�u�R�/�-2\�㋂<{��� z�X�<6�x��?x{�1N���/�-R�бq���l����V�?�����Ҷ/�E{u���ν�2�m������N-�R�e��S`a4�3NU1�l'��?�#KB�J�>�s.,�è���\�����Y������U���Q��4��h0�h��W z0S+�v=,�"��l����j�$����3C��N�D�)<)W�?2N��ZE���Z�pQ8ޛ�EΆb��́,E�����Y߆��F�E��\�����<u�yIР�1 ��{ɨ��|[�ˊ;�PFcԵ�� ��FSa�)�KG��J'e�]V�4�;�3��*��c�G�9&�N�V�(�-uٷ�Z�Y�JC:G�K�&ކ�Ǎ!$"ٮr�*=,���F�+���oL��iJ���o���mS0B����	�B���k�e�$����xd06�F�<���/�5"$��u��4�d���|B|JU��7"�
O �-�%�WǾ�����H&��q*�g/%�دx?��,��^n�c`L��e��"̆LB0?mG~��o"��L���OvL���&�8w�%���Tk�)1�D�D=�Z����-i��ڤ#��-��� *T�C_Ѐ��.b�\�c<���M9���<��r�v+��:�g�~}��#�ޯ��	��G�R�U���Ȍ~���sa�f`��4��t��I�8�:�k����b��/�&��S�S$�v_Ԭ�M��F'|nKh��+��?}L/[�x�����]�&��!�ҡ�i�����a-�&�[\;����ֱ���	]�7`x�3-��ư�
�ڙK�U�c+�$GAc5N�&���m�:��#`��)�$�4^�sTy�3��эP)g��>��t�bZ�^ח|`�֐C��H6�tz��&9D����;��=ɫԛ�Q��� ��'Uc}5Y\�I����g����Pre���fKɞĹ.Y ]�B �o�I��tA��EȌ&�g_HWV&�F�Y#�B���#���w�p J�˶^�i�W����Ș*�v[QKw�b���̔�F�5	��C�޾�_������<�x�@߾�|�yWa��|����,�iA�n����3T�Ĕ�Rs��V��x��+!'����d�I������7ߧmT��w�z񫧉r�$�z�2�U����Ag؍yV��nuk�4�_I`����
���܊�Z41����.�l4����g�p�v���j��M1�H-}�l��(������U����g5��wꛓ�Q�j�3�Uŭf�9��~��`��<�"�N��`�����^�=�H9�,i�v������{���j�|i�b�6�OC(��8��3a�_�M�Մ�m�̜TC���n��sY�b1�Jx�4�~�6+��������~Ьn���}���V�n ��܀�!��j�\�Q��s����1�=�~VFi��ka�<qyL|���V *f�K����r��v�uK�۹38=L;rb[�[QƺK1,?)p�I:�����V��'S9Ǝ��1eft���X���]m1��k(EVy���q�5:L��n [,]��.i/-}	V�3X�@tG����H�q���_����^��φ1��N;����C�&�|!v�|������6�y��>�Ԉ*h�Φ��*�2�+r�C���q�v�G<�-�r��K*G殲ƴ�X�R�ڈm�ٛ}�q�P���+�B�`���WD��D��sAx����G�9D@�w�,�k�ŜQf��e<�+��`�ɛ��C�E4̚e���ۢ���x\�Wʑ�9 ),��"��	�J�y�A���3<=쳼��M�E��"_0/����ŜD�M �<��VF�����W+�%!FÆy���&/T"V L�0P�
�V�+D�\r�;/�Ln���:J49鴇A4�hpL��M�,�+��ESe=�驪�\��EY���y�ł���w���� �$0?�������&`�Sq�����r���]�l�#�Y#3����TCv��+����K@U=�*g�31V&���>�t�Ur��`�������nUaƂZk��û_�H:F����T�4�;h�c��r��;%��kjlȼ$���LW�Z��n�E�Pl���.�|j�recש#O56(�븐-����#+�q�ڨƑ�j�� IU�����9��\�ٓ�B�D
�)��^ !���T�RԶB��U���&�k�%TE��#}�d�0�ޚ��ǈ�"� � �g@'��~]�P��V䢀����;������:�$x�X�WG�g7�ھ%p���t�*1�%H$`�]�,�k�����J+������#y����8�=cΛxeW�(�9��%���U~�	L6���0�v��Y�W{]�o���6��r�>�k��鸶.���r��Rc�Ƅ@��l�7�yu��}�Pt�l�o
�u1P��/	�B�D�+�yNi�*�r�|���3w��˲~ee�Z	W$,��eմ��<�������K���]@d�F�ve��h�����3�O��$	�؎h��A�0�켃�a$ߌ��S�#5kޜ���^a�Rs,~���ܚ�R;t0�a�����
H�\�k��!�5&2�_Q��]J�XYH�VE�8TRԩd^�:@�9��}r��h�I��7����?5p;|<��C�A|�h�[g4���5A@|���d��f���ʿ��I\��������S�������W�Ʃ������{�Л.��O:m_3��Q)0ܓ�9����ʦ�j��{_{%��aU�	�����D�K��d��C-H��7�v	����E�Z}P1D�h��b��&�ː�E|�,{��x�fٖh���&5��S�\�'�յ��ӹ��澀 �a_Zma�D��DW��.J�*a���!�;*�L�����}_!�z��O����� =7eT���O�ߖ,�g��K]��0΋[��e=�vW�>h`��D�c6�p�w"x2�1��h�Ƚ-	d�JtaM�l4zť�'���*4���Q�����������2}%�9���~!���dMk�ͱ��Q�V�t�y�lp�Ȑ��Y�g8��E�2����9�Z��ܢ��]��m'��2~�w͜�̌�d�w�V}�Qo�2�*(����!�^�Y�E��Gؘ�i�7Ŧ��|�i�'BS�,r ǋN�m�=(��P}x~ۣꋪn`���M��ń�nKIW�0�&�	p�W����)�6̘���4���,��x᨟�����v��"���͖�*��3U-��wXI9 3�A���j��X��,K��K�2�7'�H�O�����ۖ=mɰo:���ũγ���+�O�+�Jd�^��\n�Gj鐏�����o�nrc!�ܺ�hZ ����G�m��Ǯ5����1��&�	����ݴ�~Lfm��� 5�9Ͱ�����'b��2����r?�֋��.� Zi`q�F?X��_/�� :G���?n����w�E�NdHQ
~��jW>r�O~q�Xi�3��b��4���N�Ct�O�����4J!9p�7�n�	^G��};��v>4�_��Ӧ7�F�*�	Q�����s�Pt	����&�_�3�;���k�ƍ���d�`�qj�3��Nr��H����b#�_��I��	eE�Γ����e�hm��A(8��H��]�{�R/�9�V�Cg�cJ�%`��X���*z�$�����L�)W`�wۖ��OD�� )o�1�?4��;4���i�v�-�"A9n���$�r[f�����G�#��u��/⋇0�����
Aj7?!��>p6�a���y�Y�ɺ�`(�/b�#��Ɗv~���7�����S��_G}�׈��}\��#\c�#^
/��װ����=�����^9h�>��fT�#@T�.����fCsy%9�nZ�	��c��˼���=h@�V��"����
�f���ڙ�bm��t*���
�
�B�\Nw ��s+�k�r�]��h�H�.lF_�[��Tޭ�����L|��-�r��>]��VUDw��6��ϰ%0s5��D��ϻ�x�R��z�����D���i����~ 9n��3E�tD��+���C�EuYh�|�|��d�jp\��뷲�ʸ���҃qh~���S�ێ�6�j�D����5�<��Ȫ	ym��~.��e�W��2_��jo���<�5��i�s#��K��W`�Q��Kf���#�����i�trM�R޺�s��]�t�!.\��4�Q�H�s�������J]#y���{��	Z��R������[GW�#�NΫ�#�
W�����q�IM�T�)�6��zi��!�j�މ@*>+�o<�|Xy��)e|mN$S7����D){�A��)�9kn���SZ� ���5e���{�?��izGtvZ�q�B��b�w箎ۅ��ü�?�	�o�!r���_�:e�}����p�0|��o,��Z�N��5��aqֹ%
�N�4|���3o#-"?b^�A�ڵϸ�p���$*�~q#�T��FT=W[�`���'5_�����6�.�ܖ��!�.��Ȼ�GT�-�����Y�x-7m��<�" p�'���)����
<~���]/ݠ�p�W�G_G[w���U;�6���RUYʪ���d��E����:�1����m[�6��;��|=�d�{ESE�|��97��`4�����������?s�u�I�h��I&��k�,5��	�p>	,��PA�a�g%^�xj�5qT��`<��@[0�/�`A���"Q<�z(�5�U��d�������K��21���:
�Ax���Bʏ��e�䲶$�6�n�4�4N%\*(�h�,�`��lQ���`PDT���2Ո�?�;NR>�����=z����M�l�ѧ���+EK�g���@Bwن*�#k�m(\����{�����{�N�d���s�α��N}i���	��C����{�t��R����
d�>���7#��8K`j���U��o����&C��7�Y���B;��B�֡پ���c�DM�%�����՘D��3�I��g�C���e(�0�c>�ڒ) �=�SMx$�i<�=x��-��v?���q�((x&������:�1�4g�ׅ�4���q���bbD4q�enD������SW
��a�!Z7�2ڃR��J}���B(B��H�G|Q��N��x��i�C�-�����i(#��R�u$�w�`Rr�L��:���RQE���#�9�����[�ڏx�F#�.}p�ل1���p���n�k���lČ_G��4�;��Zg��5���1�ռ��:�B����!���@,{0;7�d��sm�Y��=�r�997V��p���8�RH�9���%8�9D�T-gf�$d���u����4�; ��:v`���^G*ЉJB�?����u�mk�{i� ����no�;f�\~p��+g����0��.S�6Ť4��l��T�,t{5X��W��:-�*��QDs���jQ����ќ<H&۪����-@�v��'�¢�Z��c5N��ں����q�/�S�
��u���찖�o�z�jP�M	H�����%��%~��-���]�-�˫R�K��P�'�����B�붂<�\�;,I��xN�F9�S��l@��Rm@��C���c 0;@�Y�Kr����J���!1TD\E���E�� J��Oz���tù.�X7Ӹ�|�'�z/��I��E����v}�9��D�Zq�����33oS]�)��D��cu�v�l�:S��/_i9Ez�P=#��j��W&@�\�8d駳/��;7�@�ۙ���g�M���v��ԯ�F��3�X1�Qu�G��봒�Y,�%&W.�Đ!��z�jM�Zt���~�O�mc�ن�vJ���z��OW�-�>�/8$p��|�ș"Ѻ6�ô1)RƂi��Ч��0�{Q;o���h�qg�/
�LMg���@�"Ѐ��aC#R���P�<�f�1�h	��v�g�La~�ɓ2��~���g�У�7,�m`�n��p�܌���4������`�-UJ��N��sM�* �l:(������gO	��ρ�_�^m����%:��<�V1�a�G˱�}7\��_�W2p��x�v{��tO]_�,�З���S�#z�[����n�0��#]z�o�{�WV���2*���oƕL'��#��d��`L�����E����#j�Ӱ�:x���ɟ�r��5���@$'M����}�K�Y��@�!捻]��\[�'g�6�Ge珡G����N�k��VóL��:|����'A6���HK��E�#����2���V�k0�;Њf���(]�C>	��D�����O����?>��£��f5j#��	%U������BG�=�麗6��WSݫ��%�"�|��]W5JH.O����KB��X�l�;G��q�.妀^ڮ�0�x|�GV���Z�s���g��К��_�!V�A��VV�Y���?U�� �d��h4��`K#�+n�M�����~9-�v��+�����k
�����ti��z�?��󰋀\<��c%�������T�+��o�wf�
0��eJ�.�i��yvP�R4�('�6˳�I�����6,ώ��4\�f��,���Ma��Vk�+�ul?������C�K�,�jc�T��M#��`NP��/O���7_Bɳ'��
����?:�@ ��ww�Y�7ܫl��=}��V���%���ځn��CuXH�B\��X����a�(�M�upF����a�Z�(�N꼝&a�`�y�A�}3����Q�]W#��Q7�vc�k� �'{:�k�<<�|�� ��ͭ�g�Rk�b�qR.A�l���ʌ��W�c��IjwN�WȠD<��'W�("UfO^��M'Xj9��R�T�l��# ŉ5�i/�ᙣ����� ��#�� �qLW�Y��V`@����P8;�����o(�Q_�6"&�X�g?�Y��\���y��To%�a	c�O�F+���M�!f�.�%c� <3�0 U&�^�=��a����Ё9���qS`���s,�`�.т�i�ɃU�r	��q�(#��$�q���!	�}�8+���?e����Z�.p9�����r����~�*����d��/Ì��֍�� g��\jv>�[ L-ݖ�Ӣ�@͚��)60����k���v�3���K|f�ڜ�(q�,��D�Bg|�;��t�������j��d��
"���n<xg,�Ls����HR?��(�=-f]�Ǆ��Ie����q㱥q��z�aI+	M^�'>%tO��=��)տ_���$�-Ĥ�:o��6���Ae��
�B�K �\��f��.Ͻ���KfVwd��E,�tT�M��4�b��H�iB�P��S\�uҴN6���R���B˒�-A+�kOc
I�L�AT��a�|Dy�"k���yk\4U��ҫ�m͝D�a�{[+bҧͫ+�[�#e郷O@��L�gZ���"ߞ�Y1q�^���%ن),�bNYt�ّx���ܞ�+���Ĳ�,'¦&�Iⶖ�\i�	��d%W%�E}�#������mU7�F"c#lۺ���Xr��e��;���?����V{�-�ן�p�I���zχ�~i@�~���w��Kĥ""���>s
�-��Ϳ�eM���(�Gy8@�Vq�ﱠ9�ʝ���Z]D]���υ�_M���kN3��3�o\p��<o��?�g�a\�@lV��j��\]�C=���D�:S���7���f-( xc%X���g��R���%����ts�fk���\�jn�=��w��JN�$_.%O��H�-�I�t��RƮ�q Ծ
���f�x�&L�0�yX~��v^���cý0����D��}�xS�wTAP6��T �����^�E{������5����AB������QM�M�j�uZ�j|UCP��ǳ���c�l]�q���xUc�M��z�Ld�PO���pL>�'^��@J�[��W_��ݏ�X-������
ä��<�9�]|���g7��4�a�LY`?�~��,V>��JQy]L |¬�� ��<4S(:�vb�%�� 	M�
�[�p?��&��ˡH��p�g��9��d���}r>��C-6%�`�%[�����Წutv�����T�2�Ç.��&c�C�U=�t��G}�c�P��\��B�q��� ��4.���+�gcG[K�6WS��UJ����r��~��f�\[u�YpA�	�r���w�)%�t��3��W�m���˞����R�s�!���{��|<F��.E�os�A+�6���@�\v\*�m�-8S�?�.�G�fX�ķJ��K�Q7;O�g�z�I�_���L�b�*��#cϨ�A�v0��ao�*�j
�B@tj������*��=���ҕ �HA�����z ��̎��TU���Q�3sk��-��+	j~�1y��5:/�_��(�=G�=��,Ч� y-қ~'���,E��㪳ZF�VC�Џ���?��sj����2�6.T�Ts�\(�J#R�ݏ�����Oi��3��vz}������1�J8�t���M�K�f�=bavX`b�T���]�-M��p�>+b�P��h�NH�OuT"� �,����C�����H��
�)( {2�<��;��4��,��c܃u�z�����0��%�� eR���� .��C���9C՚��R�R�=O��x��)�$��Z�|���O#W;��y���Pi�[�#	t��Z�7ϚAS�|=��@����#��vPg�^��O�w$����ˤX�������7L;�������w�cާ<�����*��޹�~@A�.Ml�Q�9Q�7�ޞAG~V+��+�QZr�-���N�@P�3�@K��Ғ1빜������}0�rJF�S�� w�������J��\ �a�?�Eez��k���-��g�)� k���N���c��!y�<$�`�O]�W�������h��Ξ�3Sk+��"eW,��4lY"(nϿ5���.�W�o�Z��;�>m�My�].oǨ���� �ob֞N�i�̈��-�1��S�y(?��Q�&�-��䒷v�,�zXCW#C�1e�ċ��;�����j�56�:.	�u*&�<}�~�D�%e�&��V����������~��C�x�w�H�I�u�%ZNA��^V8��rĸ��A�W0z�b�т���%��/a��{��&A	�q��DǍ��d�i��^șY�m"��jF�+y��������r�΁ܚ���	G�g}ŧSs�ol��Ox�������j΅$eN�HJE�+J�v�(2?��Z��������ƽedh��g(zP2����Z���r��0Hx.��w�����4�E�6�VNv�O�+�bpj��l܏M'��RNإ��6�o�+��9�s���93��%̝�fu�y�Gb����O�>�W[�S�*��؝��H#gw�����-�V-����0=��|1!�� ��r�+_Ѿ�XAc�JW�	sVV!�@{��p�i���8X��)]ؠ-��`��>���o;�c y�@`tt����M�a�5�q���e���@�jO�R��Z�#��S"�l;|x����,����2�ܘ���Y�Ԅ��Ɵ<ց	3�6�*�^Xƾb�u�@	�YI��jk�wf�X�.�	f �<����N�\�EM�Lv��kKR<�\_����d� ����UF�0r��=�Q3�{�V[=IRks�����U}���X��H��*.��(��fx,&2X*5�7�G�����]�{��e�"F�D��M��� ����H�\ǣ��n'�a[� �ado�;�64�;��l��>y�g2�
	lywOv�����l��C��ǯգ񯜼��X[�w�>�$D�d�J��X:�2r��$}k��f��p��C����*�f��Qɞ'��W�����KzSS\�6��>�En�y�j�F�P��_73� ���#�2R�9�{S��CEo��;���?�����!���'�Y�p�:6v=�R��-�1M"߰�ta-���_�"��T]L�.kV�e�A���9՘[ ��P��%W��
��8;@��."����D8z�[2����a=�1vq�`w�"��#���|���;�K�v�>�������K<w2e1�_Q�R��oNUT>�:����Zȳ^'�ěĬPNI��42��t����&�F�� -��e�� ��=���]m�P�����1�o͐5��0�	p-m14�2�G���[�9\�����D �\io��#T	O���o;��;����<�8 �lu8�_U�L�ARGÚ��NL���YaJ�[�ר���е[���@�ٷL��tʜʼ��ǡ+R��1�F�S� :�˿񵘌A���;RC`�7���C]<o=��	�"��W�\ϗ���@E��m<�;#��"� �9�b�������£ؽ��Kd[� ��M�m�6��`=��ϜU"<x��
����"Ƴ�͘^���ͼ�f���$����e��T�ݝq�����1\��	�:��i������r���O���ӎ��3>m����Xu^*��!^��^�Ih��@<��Ω>�W^��ۓx��z�}4�O˨i���r����P�cCٽ�s�1�/␔�D/��~uˑ ���A4m��	y��w�X,�s,�^t�� �Am�I�`RɨՑ8����[u�$��2f�����59 �@�9(�3������0���c"��#����l	zF�:E1χg��ؐ��neT�W�P{��4vCѕϫ[�j�>�	�h$l�JWr�*�<Ff;,2%�}�W���R�թ���"������
Ę��|+!��ѳ�+�Ͼ�I�'�}�f���Z�+6����z$���C���`�jxx�|�e����m8���H�ݎ3��;pa`��ŏL��c�����/n�wF�18�Q����B�=��'	���t)����#� M��H3�srݵ����Ĺ���,�r�9E\5�4�4��Q�6T�}���1����仑��ժ,\��/��ek�
�q��]�M-3�6��*�p~�����>�7Nn��Ct��7ϐŁ@�iG��tg�O���G ���;�p�E.����ð$��Y�p��M�O�D�O#��0����Xm���Z}U���S�ƣ�/�����!��B|D��O��A�c��6gu��q.��#�p��j��(8ξ8-R�Z~���{`G���I����D����k^��}x�i{�sb&i���#n�|�"W�ϲ��sÇ����V$Q�-���raH)��W\�)Yd�R�TmI�;�\�_!���O��챈��LGc;�g�L��8�3��N�<1Vc�Nn��I����,�D�~��2
ԓ&j\O�)������N��d����P9�#.4�jү�u�Y�M@K�Ҁ�[J��rBX�{M�gt���$�$�������U��9������U���ARq�@
��.	A<ê�E}z�қ�je��Q�.Y��i�v\c�-|��hl)�c�{/'���\K��YӉ��Sն[���4_��	\+�`�ms#P%��Z�P`{�#Tur:�P���zo;�O�	�������!�=�0�W��½]��FE�S���ۥ����
��Xwf��G�?�L�]���Wf��ACz�����FѰw+?"��78���7�e�W�%"�)�ȕ,tY$�<i1�-��=x�[s���'C�lG�'y��\*Z�7����)}t�xV�������*�r���j�:s#��V��t8��!Չ��G�:�8�8e���1p�]�-��mm�"{��-O�|UM���x�z�v〬$4,^�{.Ք4��� ��Hu���U5"�xX�(��� z�x�Ru��ؐk��W����"t1}&A��jrZ�>N��3����D?�Ș�;�	5?q�h���C$����Ww���wf1ek�?3��p�B�9^	U��xu;�~w
N��W��I*ajcr�;_�K���9�]�E%�x	�?8���
�1�$_јD94���U?��jQ�ǥĴ/7�C��5#/7��*�))Ɖ萁�>�إ�K����_����[�1�޺B��X2� �j~����̲����_���2���]A�]m����B��YĄ��6�>� U'%�зw�ܺm�����Uf�7�+������'?��=�GR���1O<��u|:dϱO_v�Ur�.�����ϛ@�:b�!� V�׿jGe�������T�s�o�<v��}�_�'Brg;�^[�ջ�������N��Z�Jb��v`��b�l=̽�-�\8�_�p�D-���Mlը-=4�*�D4���wO �%��|�N*�:�-�[� ���p�{��{x�U�O��5��7�]��ڥ��?>k�Y��3����_j�G�uJ5�p\������M�d<k�
�~�f�S�sn�~E����������\;=q����3pN~p��'GP�����o$��)�xY��r~:q�-�V
,��k4�`ǖ���No?�4�n�����.��ZN''��J�XǤ�$�Y��v.�_�<��y���׹����-�)wy~�Zj���i%ǬG�<L`'����3�ha}X{�����㯹ڝ���(���I�����3���#��xɳ������*nG���v��k��R��b��ó}�M��N�v�NjHp}n��Ű^�W�`u)�؎ϭz�=��f��6!6����A����Қ
 eN��O���`��C��̥9�߬����X��ͨ�\���U�Q��v��/MtQ/id��g.|��A@�`���S�_�i�bC���f��p�?*�h���>�-Ppk �F�X(ua��H^1����k��W��~_���˟�rR�E��� |,��q1�!Ĥq�zv�[�>�uD�g�QE��Wpe�`����y�[�0v�$i�*�d�����H���t�Ӹ���r�����n���wSǡ0�h5��f�b[2{�*,��_m�=�wټ��ehl�k�!糲�:8�ʼ��A�>\�=�oX��g��Sҧ4�~�a�����3��[��)�/h->�� E�:�"�ѡa~�>��}@�mp*r@��)Xoeh��^[Rw��Fֶ|����4�j��z&������ˌJ�G�238o;Y��V[����੧�:��B�8��������bY����у�%|�G�>��緼/�5T�%�؄�:-砆9�0��5���hE��W�!��#O�>��~1i���c��{%��k!�8 ˨�s����ZI�[��+��;���uw�
�BR=U{o���\(`�'w�P���Kb��[�2h��\W���);�Y�m{a� 1�d��u��~y8�$��y
?�F�� � Bg�_����r��`p�j�A�i���8�2��(X�6,�,�Ca����i��L�Tҷ��hS�ln�O;L�*����UǬ�Ęs���$�w`	�������X�����h[�oH!!��?h��F�G4�g��8�]�Ju�!���}_V��Fa�y�K~Q:�d�HR<[��w���#�V�uqi;y]�m���9�8e�+��k�c��n���#W���eK��`���h�uo��u���VV�W���%$D���f��S�e�bF#:�F�bd����<8/����8��&�s6�F��C���.�S�^.�o%i�C%+�/����?����Q���w�=٫�k^'�K���~E~�ak�����,7CU��]��%�c��\߁3�%�^B��k�B��xݻ�������t"Mr�ёs�1�ڛ��h���qw�n��qT�R
�!fkD���>g��v˭����ݙLSh�d�_\�͠L9�����2��M~P��d�I��^��f�#�[���Y�}+V7�9���U�3I���s��Z���� e$�Ƅ#{ԨR�4�^tF������{�u�$�W�;O����3�������@h
�&� ;�plUٛV'��U���	L��g�B�I�g��<�du���7�����ZAL��F���;1��N�-qí3� _���`E��F�9(�j8YSq!�1�g�u�<��l��ۅ:��	�
o,��m+&�Dvźg� �;@���L�+���σ�O�ꑣ�������e}��S��������<uHh����OBR.O��-=��I��p7�Lfz��'��;�&*�UȒ~���%�4�q��7���`�L��B�����>L�┏��B��>�M���޿�8��aÜ���&1$V&�v$2@1�ݟ��<o��G�L ��_F�,N���Uy�(d�A���$�<1�b��} �ـ�!NlT}�KS�yn�<g 4j�e����QL$��`�N?��mc��.OQvLz�2�3�5J��f�+��<�W�݆6�ٿ�8!(p����:e#��=ɱ��I�)�]�����*�4-d)O~^Z�:Z�ѳDFb�x�M�w)����;�� �p��/�����H׭F�P2��%���-�t<�'L�)}�A���T�m���#��`���T5)з^��<�mwK����_�-��\\���OC�,�TOv��pPt��Q�=ے�ڭ\�����E��|"�!��I�Y�O��1.7���˖}o���b+8^�	(ѱ���t��7^��$z⃄�T~D��gV;l��!�|oG��!ݨӁ�ҋ�Z��I�q{�"���Ү�	v�xt$�d|�XB�r|m":�@~4�Ns8��:��w��=����%$=���� �O�,��2�]j	����x(d9�?��B���dI���" { #V�����/�Ũ'��3�$��!�1<]��$O�_�.�������q>c�kPԃ��.�^y@d���֑�:�
��GH���ʺ�
m�}��r��b�r)���@���������@��b��۫Э�Q��ɤ��[���@��ʡ]n��3Z�cQ��P��lgk�������dx�W�"�c��*��4~� ��U@w���P�Ɠ!���G�;��mj�H��g28-���\��>FK�%c;�e��4䀜�p$ݦ���gt㓍��/� �D)��(��S�/�0��a�>P���"�w���QFX���y�q��;����U]`	��5�Y�UR��|S�I2y/�f�G&��`���k��{��{eKֶRž٣�[X��w�4׬��Y�@��E�&�n|w�#{d&��$"���8Ӫ�M���� �J����Ѻ�b$#_8ǵ߰�<���z�0�J@�R���(������ǁu��)kOU[��K�d8���5p��;�L	��e���;�\"͘��i�L�F�8"H}$,1zOfI�EL�'6�;��sExIO��d�Qt�5�}	[��x���)i���G��Ų.�Xۑ���A�l��Ce����[	�t��%U_������Bl���N �=?fN*�yi]$����Y;�ҝ�Ȁo
κtk�^�%��&I�	1FS�ڪҶ��/(���B&BķWȎTș'c7"�8��r������)�1G	�ĩH�,>�0a�<)�9��y��g� SD7��4H�2�"ȶ�[W���O0���ݔ��$XD_�����T+l�.���" |t�6�
��P�g+m�]$$�CWH���Q(f,쳳ϙ��K0w��ҠC�7����(� ��3!o�}�e3/��.ƻç%�s���^�LH��ZցxJ��?�iga���k�"��f}�����,�E�kbPӥ�;����;_�
9%�ś{&��CtQ+�ག�K��������+�_���:-�:'�yL%ʈ���2��J�t������eV��
v�V��:ñ)���r
�{ӂI�F^?����}�sO8����`���g0x�S�U��u@��X�6�L�V�RgҚ�st�G�T���AZ~Y���5?�- ]e�.��*�"G��(�"�F���!���ī���ʀ�^*�}��)6�>���V��.�'iN�A��G �a��J�
ӛV�/K�$d%��`"'��	G���c$f_�������I^�W!ܷh�U�0M�&o�)�u�|�r���q��疌��!?bO��v�4Y?6��7Lj�%MMHuO�D$��Wl��{7�<"�&ᶖb4]d��W�6�-����[2�����ylI5�s�P��U�2�����*���	L\\�Q��z��p��D7n��^�0���g/��]Ë
�\�~��Nm��(�8�EB���������m���`�fSx\_[xOL_n�x��DP���E|A���X��szo�X�CZ����P#a�N���O�h�P���\���^����u��ߚ�4?ɺ>��y�*9���-Y��
��6c8sl=�W���)��qfns�1uJ��ƌ���f���J��Ͱ�S<�䊝A1�=3zod�\�I� �y�H�����Zd�)� ��-d�
�|Ǖt���=A�P��,	IB);�cabF�!�S>@(�2�]!�T˭
�h�O6�+b�>>�+Z��p���7����Z�dd0��(��}�^#	�'�2+h��vO���N�JI�)�3��&��`��b⚈�3B6��ċ.D'��Fi�CR�w�Z�}�"�����P_� N;��U8(�/6괿52���o�	�M�0����$s��"Fl8Mr�a�M΢x���Mn��0����N��E>j����p��?�9�k�>ډ%��p|����e �I�������C�|ܥᡣA���	�JA5" ��'\/T Xj��q�p��	�B��{2i*���)��[�FIU%���#�`;����c{�+���1&��go}1�mw��53I��	bUJ8!Zu��3;[�ѱ���å�� N����/vJ�{�K��6�Q��ޱ��
Tt×��q?�sq9a�-<?y�/�!���/�t_4�,��J�Fc���%�������J�3t.��/�����Qk�5��E��,�lUm��G�Ӗ0#��q�\)�G�Ŷ]�6�0Տ�~��P��Q#��l�S0�2#��@�o(*�G�.����$�ZǾ�����S�s+�����%+ʾq���i��Z�0wL�rt)"�[�����ȸn=Ύd��Ap�P�����
2�ؿ��h�5X��r��4^���?\;�'��Ҫ�⾉(zۚ����ۋT	��5���@�IX��"�d�M�3���P���V���;T��D�T��ܣHd�c�� ��B.�cL&L�y�@��x�Au���][ǡx���z	���"w��� �J�xr��<��{B	Q&~�	�Þ�4�!!�̄�-KM@���1��F���( hL*a<kSU(P�M�A���:��`D�"/�Z�Py!�C�mԂ LݍQH@\s��n*A���"��Ke���j�� �'��*�:�:��Mr¦�����Qn�ĈR�{�	`�?��w1��PK��!�ܧ��Ot��2#��*��2�ɢ[Q��ľ�7Н&��T����0ۣ��va	q���%6_{����yſ/^�M��e��0��q�ii$!O܌S���kV�*^q���f�)׫:���1]�K�dm��|���� ���f�I�1��N�$�}�O��6!A& ���{���4�m���΅]�R��b��C-F*�b�teB@��,��׎1G�	��$0�>S�Qq�/幽�^�M��γx�����!#:�Q�Nj0�6ф;���V��� �biܐ);�H|���.�s{�5�x�y���s��nƙ�7\e�2��k��I���q�t�T�|�=�CnC��,��p�g�2|���l�����r�;���HM˚����Ck���e�r���&^m&| ÚT3nV�#���|�FG�Z}@�*�s-Jc\*�B���� ���'�?$$��	�h{��+�E0�h��A��a�7�I���S<�+:X�TtjBڡCE��s��}��sّ'�"�k�V0�]Ζ�vb?Aj��dĈ8�׷ %���̺���贱%s�k�`�_ә�8{P!�$\��i�I򪻬&&�&eg�A�9����qgq����F�[T�,g��cjr5(��Vd�y�ælY)0�p�)��8éU����ZJ�T����Z������C��f��������N�%n�V/�X�bƴ�p�D����^��`��]�&��1��*��@����>�>���ji��+g�@�d�\������/
O�C�:??ū�U+�4w��qb�o"?�P��me�������#���̐�4��Q�K�B~VW3"�(y��=A��dV"�G���K�����&*[�����8�>�3"��1o�6�/p[W�41�� ��	�X���A}��!�%������No�~�Djm�>�I��
���YWj���	��ڼ�� ���Ͱ 62�x��\�ͪ���I����ֈ��32�%�	rv�RVI����s�+:�q�ڑp�����g9�/��d���8n`iVa��#<	[m5yD�=�(��r�0��^[|{o1�b�]�o���/D3�G��Kc�b!�[���6����F���bޕ�o�M�uN,j�I�1�$EJ��g-3��9�[�M��E�q���b67�9�J(5||C��#� �^�-I����i�L
.�Po�v��K�7�t(D��2җ}�^��� ��?C�E6�3��<���P�K󷗹�4�*M#�S�Z�8��g�t���R�X�!��b��cdP���/uU�a�/b�G���J�o{a�R��/�>͌)�B,ᡵ�s�mN��Y����-�m"���J��~�2bu�0	��@���Bz��{��p���$B��!&����pX��-h@����j�����s�r��l��:!d�J&;�CW�(�h+��E�Bm���L���<徝�Y{�p��w=�Kg��}ɠV���_��xaV������Q[}'������欬��*���8�뷉��A���A���M�A�v*����F����^t:G��&����2rh��$Ӽ�.]'�u�A�+�֌a"vmy�e�*\n4�������)�!�������g�O��)\���;}�=XW�����@�ٯ��W�3_b	W�.
�4�T&��/g4��sE��R�b֋���r���d�$Ј�*ê�~/ŷ�1�c~!}ܾ�R�f>G�����Z��g;�
���7�z:�|
e�o�����j+����(�X=�B�q���D��@�p���=���r7HH���pPIF�!�һgˣ�[(\_���:�9�GA�4�C��N�6̷i��ՙ����v�1��_#�Wx�����C1�q' �~'Q�O��5�r��i� ^�W�0���	ߣ1G�)���+W>?�k߿��$�n�c���jL��}[��:_��>=�&�
�n{Ŀ�El�$Va���n2��%���?a���I�3��ٵ��^7&�8)��>���~7�H�����T>����-����Χ�{��`���0������c8G��Ԑ����:�h�����ڌ��G/���?ח3�u#�yD2�_qhPaU��Vs;E/���<����_��r��v�H�/w� o6tB��
0�5��a�`�{��({;�l+prj�\����EX�~!t���_�lN��\aXrߘk���5�5�k8υ��k��?���%kG�$I^���J׫�Ș���_�Ty���;�2w��_�Ry���(�<}���K�`"�,���"v=W��������)�wP݄��J��5ܢ��cF�����d���:��I�@���"�>Ŗ	�5�z�:�+�N۹ץU���Y��j��4���=)dx�0���h��&�o��{~���`�`����.���X�����?������LFU��2��Q�ѹ�GW�,�v�zU���>۶9� ��ú"��խ�/g4 W֑=n]�&޶�6��|SzP{2��� �qC��A)s�|.�zP�85�2:cs`�\��34Q$;E��G�fOg���Ûx*u���6fz��~�V�b����䁩u�N�Ac���ɘB=%�yt�e46��r��95C:�`IeGƁ� v�Ty��Zf���Byd��;#@/��<���zA�>�s�:}������іԃF��V+�A��J�h#��G���څEAw��o�(Ue�늮W���o3� 
�K��n��A�/6@�7�f1���-�g�f��	�a��l���zs�L|�Gw�Cҳ8���E�N��@�O���~���Y�	Q�8�4�j�0���"�$#�L�5.�s�M.s��*a���>b��T�(�`_�+n��v�Io�t}�֕Ū�\Un@Z�`���yH/=�I��dQu#��u}�s�4~�W��]��"��h��Z#k#���	�o}�@�O��Q�2�;�z�S��/pA��ư��c�Ʊ��+]���w�$�)�Q�
�i��i�=�b�X�}�Y��f����1���@'R����8���f5�L�u`C0��������7о
[L�9�*�����&���j��fF��=^+s���<
��K���a}���Ebh867�� ���\̊��VWQ{*Fe1�c��XV���bd[�E��H�A�Ɛ�x���Ӆ�� �k��E���șa�np�I��}'�Z��완� jI�����P�9���3?Y������m�Ȥ��VW��>%�J(�)�Ĉd;.�J�!�j���Z�@��6��Mmh�f�y/��8�z4L:@� =�T�G�������7cHo"�k�cfgdC/3�yu����;�E�\�5�Rv���8���|��a�E���R-He����Q�Q�
yU�h�b�*�aB��r�@�niy_TVH�V�+����^�������x� ���t7�Q�Fb�%�!˲����G�9�B��EGJd�8g�����Ƥ`.bkځ�m��X��R|��\�"���4����B�v��'X��$�_i.��t�:�J���F���y�V*��s�c�Ì4e;�Q�~Bc�u�>=� k{%P��pܹ\]_��#�d�Y�$1C�ś!|�����З���`Z����շ���)�]��^<�>�p�0��W�ͭ�%�%'70p%��v���}��,���g�i�-��
$���g��8Ȁ.�O7����d�/��va �t�ػHXsݿ��m�EfR�C��#m��dU5��~Y�+RC�W�y�ӝ �A�E�[3o��&���G5Z�H�eT�Q٬�YV+�Y]N��db,s����q4+�o�Hn��A]�v�N��e0c�ɏc���p#��D(#���>�������K�rPf�E��)GM�6VS�����m����$R+0V�z|�����R0� ��'SZ����������'9�͑�M5��ܾKp�~�%iop�e��\}�m��6�b ������� 9�>�'�|s쩑,��+ ]9A7�O9����_pc6���X�O�#��c �|��;ܸ7���Rd>EEw*_@�(���|��ha�'�q�S G���7��K}�f��!���^+O'�H�����E����E����kVƓ�yn}��]�u��xd5H4�����ݏ�i��IwNb�~���{��
�0����4�)d�ԾA Yd�X�FG��j=��b++2�0-���	�BHPi�n��h�� �Y��y臅$<��nS������Pƪ��`�}2��(�n�#�ٖ8;)������wxY��Y�sΈ3j�E����b�F�)�8I���X�yq�����H���qg�G;�q��xt�A�q� <}y�H�U�g<ڐ�e~�n�,b�Obt����䌂B�S��8#����.���(Gh8��@B��;r�lS}�Oh����S�s�[/7���k]���l�{����V�X���9�?|���>ª#�h�1��<3�}ǚ����O����FL�{�)rp^�s�Z���Uң^���;l[_�˹	��߉���'C	��4�^P搹��ɐ ��M�������!8s0�Ca�		O���!���3=ӊA�A���.R g�*��~z��*��8c¬c t�^�K��t(%����K����rV���v��&�e�,������	��`����y����"\�*e�c�.���f{7�𭥰��E��5���.SZ�l�˖��#��?����ʩ7q�1H�WP:'��h��wJ�!��}��F�.�`_�����C�6a�+.�E�8�eu`����Ie��]#���s����^� ���{5���$&i/�,9h�m��'f6*$��i��`��z"���!�g0��,�IM�o��_$۵B̻/��{k!����� �o%Ӎ̘����ԂkA �r�
&�P�����r�8'�R5�b7� �(����%��޳X�M��Bڎ/�qKye���'E�.��Q,�뭫q��"�-QX�^)�Æ}�졳K&�)I�Ȼ׸rP��6r�)_�9�60�'u=u�o�e�Ƴ�7�	��] ���!��R���o��j6,u�u��5�_�I��g11�TK�%	��ٿ��v��)�	c�dv�6���Z�448��6,e"���n�{�pk�r�T���C�=\�6�M���&D��{lR1��s���Z`)��(�q^�h�im��݂0"��ݶ�F��z{!;�jW���1ST �O�ʮ���� #����+���I�M�[^��pI��a�Vn�;D��#�����)���TF�ɫӧR���@��F�W?�7x�䥶���A���_A4=n(m��T~f��Um��CLb |ٍ�M�Q��}>��6g��T��7��ap\0�t��q�r��KѠz$�4���:n�/���p�|D>Қ����U@'�v�r��O���8�C]���Y2Y��BD���������($�G�M��Q���w>�^)�y��'��"R��M���t���ҭ&2ݽ��� �T�l|X��E�'I:�Q�L�}��Yr���@+z�$���mx��B���ˠ*��5��)�.���"��6��6P�3��p�+��oV,�ô��S����́u���KqG㡏N��J��n�0ro��텙X�3&\��ȓ"�b�#`u�=��v�Z����?�OmҟƳ�yǇ�L��dC���Y'xsY�Iך�r�4�N��	�Z�A`�;��Z���f^�/eE��W�q�=�)�.��W�ڦv��=����M9"�6sW�&���X��o܃A�ѱ�^Img�õL'�mP�T�����{�]��;%���x巐�<QI;���r�RD��Y�8�j-��c�]�����WS4Ԓ�E�g+�H�bE#��)���*2Ul�
�!�(��i��~�>��ts�g����^���<|`v��b"n(��g)�#��+���z�G����)����FK�c"r�Q.d[���(M�b��9K��ŕ:�S�;�J��O�!�8��[�:��TS����Q��$"��a_�y�H#�W���Vk�s��񖛂��M����A��-�t�����4�����y�pQ�5c$��l�{����Z��/GH��+u><����� �㟇���;뢖S�M���*�8�ZA��,w].p��Ӹ2���{�W?�}Me�m�
�6��G���8né�K#��b�p�c>i<0��O�����?ǹ_b�<2`�@�	q�U����M�@�u��i�޽S��P4��W)���K$��w'{d?�HB�!WeQ��5�hCT������N�.TS$2��
B���Cy�lZ�"�����@�}$���X�@
�Y-�Ju��\��IeȻ� �TF�������נ��&f��3ޱ�:�t�K�<S�Xy2�%C �;Ty���OI�E���\!�R��X/oB�Z%?��
O�|��d�!>����a9�h3OJ'���$>�9��
	洦��9;��&�����;��g��Fs���d���s����=�k��+�	ys<��_VY/�0���q����,� �ľJ�*8�ű6uŪ���#׶��u��G(�,9���^���(�)� �^��T�m0:/�Ɋ6uՂ2��b�%�`/9x;���տ�<m�gx���:*�A�e$r�Y�A�o�\Ti��}�����ʛ�L7�MA�
��5�ȲtA6��'�u��3��y�����eY��<ڐ��t���<y-�ئ!ԅkmiC�ZʳWɭxN��"�JٷHd,R����0���� �vA?M"1S���� �{��(��"�v�(Ć�N���̉�4��Ȼ�S-gi�����%)-,����/��/#$���N�>H��ܐV�s�=*����+Z$��D7�1>㐘-y���M�DI�G|�0��>����e�h�U�5�	�_�F����R����������qŁR�y�#n̘p���Q��?���
�JY����9c>�=�������H�m�7JW�f;h_r���,#�wC����hd�x�eb�Q�=eU^KϷ�a#2�b�E,�����-4ͣϤ�q���c���O8�
 *��Vת@�*�:��TL�N�V��JL�� �|���(j �G�'Ѐ���djjtx��)�8��5��7g�:�ֈ�)��dx�����+��z߆T����6����#�����h�Α�>m�|�"�'��7�U��FO����pB	o�JeU"�m�C2�E3�13)��B�1�~ ��3�>9p+���UY��2�	tV2`o�e����C����I7;��Y��<އ
VE���e*Ю��[�<�E��oC~�ES�/6Z陷�3�tB3����ͪ
/����7}�-���7���[CG�h˯||��r��>!��+�㶪֋�ŒɅ;cK*\���U�����2��;J���;�+D�Ҵ�
ZǃG��?�R@XΌ��\��meo�X�"�*�bU�S!em6<K��0?��s�b�Ld���1��p���W���9c�2s�B�;�e!�������#��%��v:�/�͔�Hzى��Q�/���=䋭<b�P���0Os�Z�A
ȟ*��>3���==���J��V�IU?U�{�19����g��'�d�׆S"46��ӛ�4���4?2�b����C�4'U��PN�W[��X���%d��ֲ��i]�%o`��3�������؂�}���ÓH��	�S��7V%`0��^P+g���Y49
�Z��������{.��b{�m��P'�Ș�.��M��f���J~*m̠-g�#u�nv�w+�!a�d�v[V��79���M%�gPP��$��,�r 6�h�b����"�ͼ<�̞���iZ�;q���LoO,lzC�����I�|����vks���p��b@��R�j[B�^���[�s��R��9�������P����=���1П�,T�"֘b3����C�gb�yT�W��o�.��+�l��5W$������bԻ#�>����!IVh��,��(~�gw/�¤*^�?�V^�Yܬ�!�&;�,`��H�TjI�gS;�O�V1�"t��:��/!C��ȇ.��h��j%(��������R��CU�6�3gWւ4xsL��{��"?���U!���L7j|3>���\᧑{�"���� 4� c�&�ǝS�#���N	i����7:�Ȍk��$�I�mwL{�4$=d3�$������#;�Z ��_�2K��Z��貳�9�"������VwӑA�75K ����l�4��	��!�4{N��웩��+\y�D��S2��Q�?O��[D�W���8���2�i�O��g6uJ@�Xr�'��)a���}LN����m�9}�6��H��1q�b�~B����ZЅ�bNW�q۽4x�kݸ�l+�H��f�b��ݻ����Y�x
:���z�08l��=��/�U����L�~}_���t�BS�ToP	�W��Ws����۽�\��q��}�J �W�Oo�ul�8�y�k��=u���� ;HY7��}[�`q��m�{Ô��#y�q�t�}���.�,���~S�՜�P�Ó7�j%�D���5[~��]x|�A)Z�pk��5U�b��lN�i�`�z�x���z9����`�O��B݁�W�t�:���+���q� vr�R=�n�*�IP���X3�p�(���߮6 ��&���PBS�(`� ��!�bM�3�W�d��1F��e���'_�v��R��+V���F�����	kJ)�M��K�kM�h#3�3�(P��Ϙ�����1X�����bb�
*��9a��{q���]�T����k�Y��&�P���V��B�ȯ<���[L�sRLib�.]�2p�� �o��J���{'G��� ^=�����^0+z>gw)�y;׿s�<$��ԏX���!1b9x��B�nn�L�.�&F�[��^�).k�z�� #�^h�G��x������xhg�W@��(#X����%[mc�$h�]OW"�n���$Eޢ���7ț�?8����ԝ���^�����\�,N]fwn��|�6T`뼯��1~�ǲK/������r��F���mnr��O�'�V)�v����C��<�B˻Zgj��-=m�*\��'��.���D1E�tdAgX�#ڈg�d����e�Gh����kҾ^�T��y�$Ɂ�->�.��.��^<�QG�MB��]��+��mؠ8�G0u"���J�)�x��AUj��ޜ����=	|��iJ�q"4�`��QϿ�Zɐ���|I�E7�XJ���j�9Dh�]�%��ou&�`��ނ�v��� ������
S�+�h���|H��,P��*��%>Qɣ���������;�������Ł�s�2�=Y�~���tU��OUE�� �����
�r�R��*t��USy;��_P3�k��uo]�3aa��jî���u~s`���������|/k���L���e�D�92 W�������C�u�E'�?ml���e��&���[ڗ<v�Rq���_����=$3���*���O�
����JXET���T5�+����ҹ�-�'s�CO"�9]��U=px�JF�.��`n.�G}1�Gt�-��:����Z�fg���C�����s��<A��o�S8���n�/�@��W9Hن���4�vm��m=��'��'.���'�y�߲�B� Ã���N��;����E�jx��*à�i�O M�w�=�o������Z�Ɉ�SEJ�ya�����X����( @�;1�hտfE���&[N��X�}YӮ��ۆ� �"�~�����U�_3�d��q�QJ.���j�(���s҉Q��r���5��q�n���&�$�TG��}�G�$b�/�������r�ȢA���:�g5<3b^׃QqOd��J�Ԑ��J����>�w��\�V� �$�r�Pr��k_)���f��`>�LI
�-�ѯ�1Q�O��v���O&ad��b��e(�J�ud����%U���� ��u\L[���+P�A�W8�@����ϐoQKs(�!(ssU'�{��k����`瞉V���N�ߛg��4G�΋�ֻy��6E<槟���z�[+  �R�;�D���&l�GfɅgH�0ߌQ�0#���LB���H"xoF�Ŵx�r�`/%c��P�S�ߦg4H��jNY����/���K�U�5�f���!���qx��C�� ��I�ݐY��4��Ԛ�w�IN�2��b�B�UG�h�� �J(!ϒ�\�1n`�;�xG��,e^�F�Af-ro�$|D�p/l�DO��)�%��/clͼܽģ\����������Y�6N֚��q��)c�j��H���[�EۓB��G�<��k�����Y��i]��ڮ������׹��)���FDW4n)ƴ���k/M�T���R&J��̺�ǣ�.�)���t�&��}7��#ot�
Bi&�u���ys����y��(��O���b/,T��T{1r��Ungp�r�6��YU1��ĥ^�NoQk�0��������)��8j��ϑ��2�7n�&��Dv�)���V;Ǭ3=ddA\,��*�K.��%��m�r>�����|�F͓�Cg�Vǫb1��aJ���}�+��~��=CہWa�0�!'�3K��76qյ�|�[w1��)�}gaJ*\e�qu�@�I�G�09-�����k�;1�mY���.�-T��(C��O.D���djk��Q����w3�>�:�{d��`G���8ԁ��/ԅ9�-�i��c���sGTP��7A1k���M��l�I��w�w�&�c{�YY)tU�V���E7�;�;��;��r���,i�Uxj�H�3z�Lɡ���[�����P�t�ɚ��{�0l6걧��6��U�i�o �Gݱڹ4�w}ə���m�֮����L�Q� 9�>R �����[�F�z��Vg��!}���!'	d&�^(���=��י�-�me^��U���\K��d:wbI��uRt���G�gv���lt����k�#�c�Q��V먬M�)s�(�9tݤU��Ӱ(����÷��]�Z#"96����(W��NCQB����8g-�A�G��[r_�A�fg�X�H|�3�xY��s�W������Ϟ(�k�ֶj� ��%�l�`��N�Ug�J��	����)��3J��$���өl�C_Bmp�o�稜�G/x3��@W��M��=mRd�cB�ej�r��gy"���~Z�_}q(�,f��5g)y���_�G՗�6U��8�+�a���}�Q�0v?���C�x$�u�����24���CG�Ș�� �N�::nv��^���=�����V�Uc�����Uʗ8�Պ�@�U�N�7A� �/�UQ�G=MƦ�Ѩ��Q]\��w�Mv�rV�An��G���NRבMY <���3_<��gr̓�@P�k�R}�������oE������0��t~,�ϑ�<��qJx)�\/Q�7fz��	�cq�`nU��[�����+0A���0>$.#�&���:5Q�*�zs?��}nRA>�l�k4�U!��Qc5�|o�ـg��s2���g)�/wl�C�ƍ�-��V���Q�i����|I��-��S)�`ԉraF���_�P�u��41�܊�����w%CA�h���vpD4G��U0sO����?\����D�WK����h��yM�YL��VI�V����
L���~�!�ݿ�Լ����{��3q]��'���+�W�""����|�n��Q��Ai8�̇n�~�K�~d�+J�>^���s�78S���3w�k!- �z�=tx�E˙�N���2���p�G�f�y0�4�3�6���i��M|���G[��6J��}�j�D@um��0��Ğ,r�ZN�ԙ� %�|ǁ+��^Ꟶ�
���ks�S���wpMi?��/���e{�S+��P�@�kFA+������
A���ٗ�X�"��	(��g�w��3b\N���f���ǿQ� f�$v�2�+�(��Gv���쟵Zy�@�12����#�ֻ}�g���g<(�5�K�F�E��!�w幤%F���n��<>sY�_�i0��lFj�����`�Sy�?�
F��"�t\VV� ��9I1�8�g�(�J��_�9�ZI���',�H;���u�)M�
�Y��h�W�K6-L�z:y��ajx�{�P2/r��G�a1zmq8��-�o�u�4A��7�$�,u���a!lޒ�5δmS3��AMu(M�^A��`̳2���@B$�SC���9�vV"2�.	�����%�Һ����[�7�}]���I
n�X��[zq� Qj��-��I��h�~B4e�����:�A|��ޚ%��O��:�h���d�RY����V�a�o������E2c��1�E�.��М�D�f��p��G�V�g���:3Pb���Gb�i��~k_" �n�Qā����gWV'hIఽ������QN�d�J3��ګ��F8��6ʂ<hE2+͇�m �;*��8%�^��Ӊ���^]5�j�H���M.OۆP�iwn��d`���	O�zŅ����E$��_�/)��dz���I�w}���>�Ó���r^����L���?Q�2%���S���ұb�5��3�^]�3D5Ydr� .X͕v!\*Uv�z}-�y�Ժ�.Ma�>y�2E��)�>��H3���
���_�ցk��$}�*Z6�_D�:�xB�Q;�,wJ2{�4G�G�5`��'*Q�?[��K<rNV��ii�ļk�ȡ�5���;
h�	A$�'vztSX��8�GQ�Q����6��|���3���&�]E�u��P���f�]�~��.����rW�Ї�c�2g/}J$$���Џ��n8��w�
)Bay=�b$TOl��ϣ�	�a�u�EaI�*�ğ�yMf̪҂�:� O�����=!PD���v��]Z���Ƨ�:��'Tʻ�T���V�(VHjguX8��hb���Y�%$e�<,��������yt,5����^��+�B��a?dA�_-I��jH1+e��>*fE"�y�W��]x�3 q�J����p�x:��:~]��\��t�P���٥t����`L"Y@��oh4��8b�P�7w�G"]������$jk���լ�ɠ�('��{qj�0Q� :g3�zl��E���K��hf�a� ًG?BM�D���P����W$0�:<�G��i�-{X��8���
�}P���S�j^m8ٵɓ�7� ��"1NR�@�K�]	o	��&�yZ�Kq夺B��0L�d7��4O�:p��G�� ��i9Z����¹�w���ں�1��}�<���l[�sS�A3������l�Lk00y=���D �t��I�§�mO��R�<��~���·�r��L�[	p<O\�9if��[�]�(ɳ#�祸z��=���<uUGz��7 6�d����O(٣cg#4.gNH��i��2��b}5I7��!,�e#&��L Z��Ģ�e���&�����ڭ��yaԎ;��@k��Cb+X+=�z����w�#�2�O(W�"7 �)E�����,�X�?�Q,!���i��c_�jB��L����u2��o{L4X����{:�C��{�xjOk����<��Ow�'���KVe0�8�%����Բ�r��^8��e�L���XjB8h@J�(P!��������|�­2��Qe?�'[��zm�8�g�8YM./pa��G��@<�ߟ�Ͳ�H<�y+\`fU�j�S�*V�
�:$gMcL�4%|81�����b��3֮�;oB��]�� �$l�F_bey}��s�CoE��A��g>�;������#�-�2r��@&�h�#�
����6R�Ie
'�$�:�^`��G-S�u�Z��ir�4�;K�U��e�؂ڰ[���2}��(���-�L� ��d��i�ᘝ�zA����m5uMܿ/�SC��C}�a���]>���/�m���3׮�f��ա%<���A�e�fݔw���ͥ�gVr����8k��6H���v����a�6�o]��-J>��F�w5��ݒ8G����I녴�a���w�\h
E���~ي�t,����dY3�]6̵� �fr$Oۚ���b7T�_5I6��aOF��L�Z�rg�XQ��Yi�&�\�K��c]'r�u� �=�ZIrq��i�]j���'FֹP���3��b�q0��tZ�鸡ft��cNp�f�"u�J��j��J�;�Qʍ�������=@������۟����^�Ub>t���Aی�6��?ª9&�$��O- ��&T�0�L`��"��Omw���Ok=�@5MDl4�u%��C��'�5e��ăiƜ.[�ހGP_�7	@/ ��g��|Ʉ0�C!/���VRL䰴9�/�i�g��Q��f������%���P�a�`!aZ�1]Ķ��a[�y�*��X�;�I��/gM<�/oT$��C�����+t?i���̝W�i�6j�^��v4��)�r��H3��k�ϪS
py0=0	����򎙐tF��������������լSݧUV��Vz���w��6�\�"�_��ٗM1)�B�mHh�1�eE�#?�F@�?�_���2��ʘ��R`��5e����I-*0?k�sȞET��A�s��ur�  6�o��{��F��;��G�y8�T�N�1�{>#�_%�d̅͌����ݼ{��t�m�O�.�		fG0�����@��@�5m�dB�Y�m����O�s`jq�<�����	�mo1��O�9#: {�	�Na�!��x	���Ho�5�\�\��,v/�K/~f6_��Rh$yb^��y�!-����:)I�u���Ē��З��x��gC2($ǝE٭1�sq�2��b�[}�Tp���vk`�/��{��I.����g���F7R�a�c�c�\Jf���:h-O�����t�✦9##�����w�a3�XK�{��r�t�,�'�c�nFJ�{*���f� &Z���x��Vс���L���}^b�(����
��d���څ���
Pⷧ_�\A>�\�34ƻXj��֊�b[��_��A���L(���V�����ul���#Яa0X� ����}��W]��x�l�!����Ap��Պ��CR�~P�\fY���:��\������� �8=1��!S��ޔ^�B���1�[����𣮌�a*��{tô7�I�%�ǺR�c�Dt!Թ��1�v}l4�
&�� �?��%���l{
0��q��ؒ�\՝Pvq)�!����׎m)��m�!Y�!��ȩ�ٺE�]2�ŏtT�0�WI�M^/֋����R�p$Q@���k�<��Y�����~Ÿi&��Θ�]������z�+@*�8�p:��#	�zK�˸�3cp�9q+୛u�c`�=E:O��	5�Bj����EH�-�I�&v�q�Z����R����7c$�JW��H��MV<�x�ym_ :���HNh�>/�m�66�{��w�xŐ4�ŌaIr]���X��A��rF��{FWt-1c9�<�1�07S��?��J x< o���-�coJ�)W��;Ue�OW��䙏=5�"�Еsls���e��K��F������G9�w�d�c���X徒��x����Hl��f�d5��+va�cM9ԩ��#��) |tP~��.�b�Ӯ}]��P*��a�e#F � ш��|K'��\�
d*,KS��' KDB*��
5����ۤ� D
1k���*(3��^��0��x���:$P�o��ә��z�p|���ųBЉ���86������*V����`2�٠����JM[7���DJ�E�^a3�R� >��k�^�t-}
X��
��!=�::#���9��sv�"U�Hxɗ(��9�C��E*��	m�ѕ���8n��R�4[���l�K]jw��PG�4��J��֯�PT�2r�*��@���[/���l"�X��b�-��)ؿ��61�|��g��Bi�����ex.*�����J`i��3�w{�� ��Ҙ�5���Z���8TB�4�9J�6��K��x�sːڪfԥ15�;��O�Es=:�=^di�P���z�V��&޺������bF����d�4Wm��y����"���� �O�2�l�x��]2i��Ƅ�A��f�h
c�![�E
� ��c�r��K�6.?��W2O��C.�@�M���X�0���x6�z�]���f�C��)5�/Q2�V�d|O,���8��anq���Vu���3eu���8�~Xo��5�?ߊ�-��zL��6��t`�����Ty-+�����nU�͑���������r>t�0�/Ů8��F��y�Q;8aLLy`kCP;j�3�����5�H������\���~�k�Ҙ��#M>�����\��Q���B��Ñ�_Bwr�*<���z��Q!r�Be��u�n����˷vl�3N[��+EO'�E�?���pj�.)t�#�O~�Gpq!��pP������\�IT�BCg��~@����X�"#�ݻ(�G��YY}� )���c��;YӞn/�o�X�HJ�F�l���ۘ�˫/�<�G�!>"1�����lz�Gsj�E���1S�{n_Pލ'���}�w�87n[�ϭ��$N'�sk���|�Rɴ��r�������bl�Ы2�cvEqK>g(A0�Ћx�g��8�_�/?\�U
��Ɔ[�
���s�@k*�:|�+����v<i�������_2X��)&��@!���M��z�̃&�r�%,z�y����Z�]��wh_%� H��g�'�Z9״���|T�U�,$��)��V�lQ�������YA�H�LBoȐ:�I�lNZ2��3�Յ��/�dӓ��\[;P�;���3�����沆������!�fU������#$��@�3㣽y��M�
v|XF80�.�^���`��1�t1� ����
H� wy�~ϩ�O��gB�)���3�'��P�O�/\E_b�Q�w��߳��� �9-�̨���g�m��$��(j�h�{*n����Am{�??�ۿ��X:��o75-Cc�
��;���I�>�-��՞ߦ�.��y��+W>�BL��p���_�<�sj,R,�x�4H�������JKI���1�ܿ�u�h�>�Ē�oM!�ĝ/N��KxD�
���|1�LR��v����%�$�1.�l
���䲻��!w�&�v	���"���g��1z��Q2�|��rd
8Ư� `(�Я���E���b��ޥ�N�i�v
%�sw�9XYK�W*��]l#���8C���%5YY�!sl���[~�q��b��&>�5i	z�]��?dl+̈��ڲ̮�����>Pl�-�L6����)�N���sӚ�L�
���G��Q� �R�k��a�l��19��������L}�.��n4r�C��\�����}=�Ŋ�����U�`S�k��'n�
	�iv�G)|�$E��bdڞnC� �-^7�v_�Ր��1�Ze �:N- y������x�X�U�F@s��Ha��Wf��B�c��_O�i�)</j��+��#㎠~��C��}�j[	h;�-�����\x��/�9͒=ސ��.6"�h�Ś=U�Q(~��Y�n��� � �mwQ���=@�PAr
zx�[a��hz>�8Ya����W��2
���>�YcQ=�d�,��O����ɟv�-�?�nt[�9���t����`�_�Dŧ��$�ov��T-k��|WO���� M���ӭe4��[?@@3U��i��Vֵ���
���$�u�<~�E7L�J���R�l���eٿ����Y�и��{/8}�c����7�:�����uɀ�zQ9�����ue����0����P���<����iӾ�ܭ ��9=!K���k�Y�z�ۑ���"O��'BD��Q�ۧV�C=:HL�Є6�ʃ�A0T�f�\��U``E�"骯w80"���J�B!k5w�Cc�.W´���� ��F�/�>�B��MP,�BT���6,Ù���Z�d=�����,9<y<~�Sw���vh�~Eܸp�us��Sj��k�=��[A��W���@mN�J	Z�R�v��u'���@ �U���ƐNt����uU���T`-����E���O���<q�����㽨����O��}u�G@ݕ얽����}��XpL�.���Uu���h�zc�%H��2��M?�s~��e���S."'q�Q7�i��طL�����H"E�Йsh(��ߔ�"p0�
^?��M��X�����|�wah�c�;�8�=c���5J@C�k{�h̏��K�ԕ#8��P�M��x���X�γ�;����cC�u�r?K[���>���%�3� �V~��d񹖊I�Z}�5wt�^�|�ځ�%�8������7O��0��F�n.��"�r��|(��hưQ���w�v�/���4A�>��A���t����te�dv��wbm���M	J^����G��P;]Z�/��T��0O
Ăy0�ѳO���q��/V���*V���E�ѻ�>��G̈́�T �4]&{0]!˂Kޅ"R�\��>p������SK�=n�`��19�]bʸe>$�����%v
*�����[�L��i��x۹a)Q�7dHR;W^Aă�q{O��9��*��*Iz��i~[����(2��ؙ�MVD;*����[�ydY?��Gg騹�q�H�4� ��\ 3?G5H��rƆ����#�ᜌ�&��>��.-��J��dC�N�O�'m�T�/ �wO�kn%$�Ŷ)'@M�ÿQy,�=
���g�3f0N���U�Z�e`�D����1w.���b��~̘de*WU��a��<|ث4Cp�^�������&7�����G�W������Y���Ҁb�H�;G5�03/���
�Ax���R����
�`�mC��RRS��j%� ����|�(���]��\7�K,�4%{�n|cT��Է�~���pn(���wF]��ZG��iO�C�T���ܔ4r"��k����w�^��l\��_H;2'����D2���hd�>�_��׸e��GN�Qw�yvi2�K���0�'Bb�L���b�cS϶F��"�mβ�l�&�([���k��B-QD�ۼ��O~[K��9�e�G��{E�^�̔C�t��kЏ�����a"0G��V��s���d�:�S@y���Z{};b�=}��g��$�Bټ��x�j,��c�f���z�;�?x���&���`T�껛2�@-��A5��?y�7sC���7��Z���WK��5EK<�e������Sx�e��	"�Zh���)5��`��\��j�o�E�/�]�e�DzOP���e7P��D��}q>"��y��zUeD�e?��@�o)o��1S�O,6�����s[a�]����>��(�@����+�Y����I���l����sS�.d��H���*�*q�\��xK۵~��̍{���h(v��Ȅ�--�h\�8!��?��% ���6 �г�yB2�r�=�} <M��=p][��;�'��z�ɦ�T?�	g>�A����}W�z�����Q���0��A߉+m��ZF�RH��C����,3�Q#�$.���5�R�>��2���*oR�[j!l�!���9���>��)��g��L�On:Ԙ��E#=��WԀ�r��S�����t%<ʰ	]�E3M5�������xN!e:��?��z�����< �6��N��V�l�𰬕���Y��>Z�q1����'�d֖ݗF���������I��D��ֳҳ�?�N�H|�^lj�K�p����'~^M�#낥��<�bL�E�-j�@��~F�s2� �z:]#�~i;�'Ч��g������2��-d����Q����Oh�x"��,#4OVW�4P�H�o�Z��%ѻ�B;����&q��)ѹ=aP5k�qi�Ic1A�e=1J�f�����15���9#�V�}8��V�9�L��6!,�����/9�A�!��1�tߤ����**G�"&y3�ƿ{Oy+�X�����تK/���)��䅾2�Ä�E�K�g𤒥�ы+�I�SH�>�~�R2)]�_&خ�cu�N^��#v���=�}e1̨/��~B�1��������w6Đ�^�U�s��?'����#�'i��a���ge�n�Z v2O�!�H<\�w����+��j����$a�������X `(l��:�`��� W.e�A�p��~=��������	��7��G	���ω�� Ae���_��w�\�A�1i�tHͳ[��g�٧���?�ۛ����J�e1�)`E*~ѵ#v�r��ڂH�D���&mG�����)>�5�O8���Av��)˼.v�EA����Պ�cc� �e+��ĭ@ ���Ky�7Ƹ�������X�sM"&�C.�l����	��'`�C�[��Ӂ�˄�H3�8s��8Lc�n�vy��=��]	KY�rn�gb⹋���f��+a�lA`, � �)-I�^gJ����$��kZ�oy�B��P~��h�\�+ƻ��2m��p�[�^	dAF���ij;�x��M`�%�߫��s{���:Q��^��p�
M^
X����U`5U�T]�6/��j%a���niLZ�"�>�&�7�5A�aMd2��/f�pΨ�x�,%��5�Ʀ̱~�5�я=zw�ù>�p�J�0M��C��M,�2�[ٖ����YJ���Ull��2� T��3��Ϣm�9��kX9$h�h@�f����~x�7�q�|^��s��+
��Hd�u���;��$ì�I�3'��_�4�j����b�1q���%�Z�����Ǝ�w������uz1ޖ�ȭ��%�~)������j�/ŏ9��;����+��fy����.�}W�G�ѱv�V<T��.V^4���8��_�	Fw�#8�iM4"�6�p��բ�6)����v��u�D��fI[=;N���5QJm�$��̩;���n/Q��-�P1�Q�S�^���m �x�[-��`-8��H�Q�C��B )�&���^$(�`��4�A2A� ap�XS2�ٿ�~��)^SN���BR�Ob��K�̿P�y��|��75�l�������w��`e�Tc���]��۠+�wƨ,oŞ�){0��&pEȅg�@)'4�p�k��c���b�2����Q(���t:�����Y��WMl(������z�чu�N���o�ҳ���M¸j�v.<�p��T�x�At�zT�tE��9 ���\h7�*=Чh��ZП��j.nx9�m8=ֳ�N�V�¸B�&����n�4ڝ.A=�A��2��� jƪ��GQ�0�/V �a���^�)M�ᑇhL��S$�+�M�Z+�@��L�#���KI	�&�9p��.h���������mԩrE��'�4���	�D~tiZ���G�hTx�Ľ�
��M���yB�0L膮�ԁ?F-���8T����5�Y�l�~��]S(e�OY]grUz��:P�Z����=,=���ܾ ���~p��̙��k���+:�y2��Gh�ۼzBVTQ̬r��d8�U~$n����J�9'@ eØ�<���p9�=ȓn�_�7����h\�� ��D��y���_��XN���*���kY�+[���o��[(E����HN�Zp@-�l[ykp�����<�6)����O�P5 D�w:���lͼ$ܹ��ة�3�R]����B7>���t��p����WN0.������XkG1�HC�� ��=K�[�r�,�8���pº�6MُD^]C�א^F����Ɉ�������G6��Ӣ�w?7U���#]���d"�E�َ����L3�+`��}�6�z�1���s�x�����-bĸ����V��ڈ����h���薯���-�3�Ua��n(n''�K�r�	�ҌX��ˎ�����J�XG�I8��-m��- �o�@�=�V���ˇ�����C�8��rA���a��Y�X��(غU��l��b��x��c���cztJ>gZ����`�8����r5ʩ�)\P�q��ӟKh���'��Rb��	�9�rzI�"��t��q��&�I/o��~M6�U���U%���R0���`q��&\<z銜�ܡ�E��h,Wy~�z�on,0ձc)�(����X�j@v�2��1N�"�� �&���8�:(;mZ^���m�n��v��҆�d�a���5ď�����B \����v oj��L����r��v��(�/�t}��I��\���~es��P;C> ��̺�eOߢ	��VA��tGf�Z�f�:;i�Q�SVCQ7U��BY��l<
�vik�j�^�+�ؖ*|�G��1g������DЅ�"o�.��l(���QX�';����fsޜ������C-���M��y�T���)��Q�#�������yI6�|�ad�쳛k����3�1V���V'�1�����UT�b(���� �Z��~�߰i�E�w5�);.�����/�f�,��FF� �>2Ǝ�2�?&�'>�-�<�c��u�f6NC�X%ݍ��;u���Jf����}T��Bu�x��"�(�s�����(p�";���g��֘��ۢ���j�Μ3L��*<xh8j7� �X	�A��b�EJ�	���_-�l��AV�4��_��T�|1��A�UvB�Ln�ʁ���u��æ�M9�\_��I��f�^� �Hg�)r��B��n�����@V��5�Mi��Id�P��u��w��L�b�ۈr���D��?Y)��A�jƳO{msWޕ�q�yv�!c۝[�y T^wo6��Y�o��ܵ�Y8Ǐ铲>�W PN��Eh�~�-�KâcEN�wG����+7޾�e��s	(H˚�ΕS���I0V>�Y�ʵ�/�j�$�S�}Z�Hmu�3�eӠ̕_~��]�v��&�'�W�|k��z�Wxᓓ�/�A����PJ�LJ�����߾�,f��=��"�j�^�#�ޙ����"wmP�[c1����*�b�x��G�z�3�9�'������tWxP��Z�K�4�mk>��Z+�>�yHT#	bY�x݋�2tg���io�Ha�xu�G������	��S�T ��2�-*�J>=�o�X
1oX���R�[j�ǻ%������Z6ґ�H��	�������.ݰ���c��$����s�V�Y��n�:c���?KV�8J5���-~�?&2oQzn7*χ����Nj��m0%�@
lG�u@C���V���3?F�)M�c��/O&t��W�S��S-��V7SM p��÷�tV`kA��5�@�%/��y(�c�e��%�\�!8��g;ȸ٣Z�N��إ#�P%W�q@%���ق��:����K�}@�ysh��枩��a�\�vQ�w�/�y����O�Z�B���D����oFÀ2��]=��Hlg�b����l�p��Ƚ�Q�~������VLM���L
0Q�����b�&GO�br�ʹ�L�����ٰ�ǾI���V� 4{���N��,�/�G<����*�T�܍���z���䷣6P�cO������	�������Bш�a�a3/��`*�+,�;rЕu=�rueH`�	������\�ΉF��
��դ�	29�Pi��o��71(�
�'ؠ�^��`�,�0��k�D3���J@�nAɴF���i�`<�j�m)-_�@�+�Z�_��H�<�׹]Lq�7{�g5�+�}1��O�Y'��ah)v����:�c�:l�t�C�@H���.@��M ���#�hn-�((�|_J���7X�ԡ�Y[��.���;r=���@���M��]�H��7�<N���z���S?--dt�о�#�G�SE�Q�1�-d�7\�wC:�nLs�07g��G���?w�] PR9e�֡i�o���I`��-M�)���eGr:�I�ͼ���	}Bǻ��ʐlg���:�vwc��ڄ�ړ�&��3gF�<���<sx(�
�����P,��8�۟��?���]�BWJk{A�G��찘��8�����=Ы�ZUw��OL��R[����x���+�Y���;�n�Ť0V(�WX�A��q�i��]�-�W�xʏ���v�܅5�@�- P)j�m
`a���]��蠬F�^� � ��6E<M�z�أ�?0y��"�
��c�v8�u������h;�%�����%�Rv��x��HBʯJ�.�sxl�QX���t�X�I�{�k-�P���n!3�]�p�s�A�J#=4�t�� �T�6,W՗�E!⣫l>^˚�O��(1-�wC��D�T�=1ӝ���^���Ud��ƃa�y@���,������c���)�
��Yd�$�y.�!%̸��
T�*��V�k��L�Ev�Ӎj9!)I\�m�?o��0�KZ��`�EJ����*�:��ֶ,`u��x�����x�HC*��I5X����-���dl����<�ZC�t"m�`���g*�KoƗ؍�.�W����F��c�}:�*�O�)l����{���R��9�d�N۪��̦F3C��H���]$���V �[V	Gĭ���B� �D��M�(���H�K�����?�0Q>#�Kș/'�tb���:��]�m)bخ�;�!X
�~×�o�P[�k��#��Ң�.o��.���/l5tʶRL��Yq���ki�l=-Q-�G�/_N�E�@����N�`1��{����ST܄�.��4�q[�P��1%|Q<�C[�j;iaۊX�XΘ��ʏ�g��UP_HܪȜNi�Aڼ@)��6L2ݥG
�_���1���ΛA�pʊ�@�3�3������g���; �ɇgf�o7�2X��|F���v�(���iˡ�*d��MG�1�K����8�����!��9��wA
�7��@Ҳ��s �����Y�[�/�H����xJ�	8�Ql��hZ(N�	f��F�#z�~��h�rݏ�$�o�$GgH[��L͎�C�\	F�%��RY��� �-���ݘ!f�gD��h��f:�mU���(S}���4	 `��y�|\	߀��m���d>��[�G������I AS�
�`X��qy31���)��~�ÖG����N�?�BG��ʕ���Q���Z`�Vjn��RrD.[�±e^d�^,o!{�6^�P�����Z0���8�O.�\��`y� ��;2E��
5�Lչ{5���{E��b��r2N�S�z�>E����\���ӓ��K[�0e�K�'�1Ѹj%F�\@���X9ȓ|J��φ����l��X� �u^8�M�%�ƚ���[M���X>Q<Sċ,���˯i�8u��_��R%�e�x=T���ߋIvT�XX?�`���aoR^/��ֈ���"����6�6˴�P�������yZ�&_���1�S��rJ�y�(��)S�v_��_W�����Ԉ���7ޗ��ȉ���	��e_c�W��j��<�_/��r��1�쮧��O�d�)�}�A���ė���	���{a�����T�y���;O�t(v�dpJ���"w�S����T�R�(�r�S�/��7�����D/w�� �z��!G�g��U��b8a�XY��c����{RtHP����Y�Kش�.v�

Nv�Q�b�e����RI�O��ʼ\�i_�$a�Q��+`�G��@mt� B\Z�aTzZ]�+U�I�P��0�yWȰ���E����#*2.*'F�B�xu$K�LюM��wQS�~>��L���l�����_c`\�7���MS鱧����+Xx}`h���]���ʸ�T�&����Q2	�m��*�ة�賵��H}K�\X˂<��".����Վ���6Svx�:�όF%g��; ��G#�y���e�@G+���s�|�+A�5�n�ˌ&o��ܕ���,��ٿ���@]���'�R����s�L����y���Hy�fS�is9BO���Ku���r�.O�
MZ�ɲ`�Z������<�HN�Ѭ���,,p}����r3��b��)�>�� ���N>c��=⋬����	����}����E���;�u���c�]�M��iaE2^��ѲFu�	�Iږ7��L����V`1ӺM��Oӵ�] ����
nr}�7Dy��W#��Ruo��X@���ty�/�3 ��}��X�d����n�uy���Dl��t���x�r���{�)�4Ͽ��,H9�L*k�9���H��$����SI���n�R��M�O�?`b#|�d�&/kw�wv���/w�h����E������N J6e��:?�Hl��P�V�d^,�:j�C=/�E��L��������e�o� ȼ$i�Ԃ-|����n_�#������j	�Z(+Յ����-R�8�.�L&�96����w���J3�q������=U��yud���� A%I��N���>��;��W�B�6O	������K85ekdH�Z�b���TE���*c {�� e1�`
���L�/�Xe�AJ�(�NKXz��Bj3(p�=k�D�\E޿	M(���A�9b��?�j�����oV���*O1��(�+kG냌|Ko6�
��I���`m�U�̹l��������Ŗ]2I��£P[OӴ�-v��ULm�&ze�DæЂ�Tҥ?!��LS\�9��-���$�����`M�/ �$0�}�sJ�0�^/�X���k��BP�:p�Hs�X�X����e!��V���TKr�*m��e���ˮ�Cq����T�f[�S+�_����q)|�����
B�7�w⁉UFVmq��9$[�N�lf�R��Y���]:�\�j:��{#����T�W}�������;uH�c�..�q{5��{�u�*��K�7K��Ǭ�(v��Z������Q*���חſ:��&���hqj���uzRW� q+�y�Z��!�L�����yq��<Y.��E�-��� O��sCq>�8�y�Q�ʯ&bh7A�������B�$_��s��
��M!*�B��k�Nl-k���5���7�fa!U�N�dEu�d�wo��*7�oճ9vP� W���sF����2�@C��iA�J�ȱ�ʓ	a���|5 D{����Oʐ����)�LJr��p��w�1�c�Y���K�aIH��������1MrA�A*�q�Z/$��;�L��\b5��ۨd��^���v��(��u��-.B��ADy�ӥ�M5�&C�|:���|V9�N��Ѳ�� 6��š=�M$����]�g��`g���m�CfR6��]��YB���������O�4��e(��or�;�F�hJ+�x�k}�����e�����O�*�~B�4��nX�������ᬕs�c�P^��M�(�9�Ž�������^�GP]�c�$�'�u�Up�!�PHm>3V>��s)���8�kҲ�G=�c`��ǥ|�g�$��wf���q��d�
1c��TB�[�G�TH�9я��M�Fє�A�Tz+���+�F̝i��%�x���b�} �EA��_)L��Q�Ecѭ����ûs��r���ڔ�¨魢
��_E������Vm���ڟه�����u�4L�3Y����Nݵ�G���|��|�V��X����8���b�s���W2I��.H�*��/��ض���%������!iWӯz\�)���6�.���@��s�����}�ޗ�"f$qg�|G,J	�ũ�.�7�P� c� h��i�}lP.u՟��}����"x��� ����X�c�&8Ȗ����A6�#$������f�^<#|N9��;�ZVQ^%;��J�ʇB��'��*H�����J�/�yiC�=�D�u(	"�����b���7��c�d	k�Ą�&l�!�y��]
]rG�J�%�S�Y�8�DU��� �*,U���J搜��- q���0
L��UB�4��]U�(���xs�D7\�3�<�۟WW�B >udt�_w��&���� �0��1	
�-c���Y� I��MT�;υDfw�d��Mz�yu��g��M\�ԗ#Q>�z�Q/ě(߮�l���qW���Ցm9$8��F׮���$�����>��#�'��昭��q�h�^�Flg����K�G��/���c؂��ZZ���֐��jh���H 7g���4��|���Ҏ��뢐,�^�HԐNbeLd� �-K�S4t1�����J��R�3����󇞊^�\;5#�;��@1F]k	���j f�d��φ�q�a��R�����.��?���x�r2F������2K�	&_0/X�ٮ�3���R����b�yVY�)�L;y�f;Y��],
Pv�f�?��}��OS'��F�VZo"Զ�K�Cg��<?WD(N��/qb�W�r�o�ͨ4�M�W�^�t�0	��f#L�B�6X<@�+|o0�3	����A�o��Z���5,fG[iT��H �#��A�����b���*�-�g�O�� ͬ�$���_F$9��b
��R�}����P�Ta�qoF��y.�.qC����Q�/]���13�K{�V�õ�Y��\�o:c�b;�ޖ;���v݀���ʔ��Ӧ�[����s�ȿ\h�|�!��c4�@5�p|����N��v�ó��n?�ԽP�8��r�Z�[A�.C�2��K"{ݾ@��i[R��z�E�1��[�M~��y?a�B� �j:�oT�f��J���*�:$NW�8Y;��s�F+'�q�����6�[���}�!�&��`���,�D���q���._"T�W�>p�ٷl�8�U��(���%lw��Ns��a�Pz�~-% �dï�6�[�����>ei̿�����DN�Z�Lq�3ٵ\6����X �z�����l�5�]�V.3�	��Q�j�{��nW�v�Gy}��͢y<��:���T�����Ѧ�D���؈sQ.BP�slW2��>(q���n�_�:&��y��k">�$�˃+Js�c�7w�XW(5"�)LQ��q��.- �����X���g�0�� �@�pV
>� 8�ӕ�,��R���D���ǲg�_�2p��8Q���̫B`^O����Zi���b�-��'�9&�I���.��ctW
@��}����e�(LA<L�v����T�8���Rξ�yj�}�tS�
mD�A���4o�m Xp+@����A�
$(�,�z�E��үHT�n��F舀1'��ṭuq`ap��b#ʈy]8H(NX�a�l{�s��%Y:ɑ+e3aJ�w���?�ύ��sJwƐ�y�����S�]~ѝ�9��	F~j��Jw�eA���G��D�c)�q��z�.���c�I�~����l!���ś��
���$Ah�GU�F�C�|�Â<�b}[	K�і�x2\�jU�}��)��w|��z<(�P���)=�4��F�La��)�x�)�ʂ��J�Ƕ�'Ch�ЩkO�l��1��z�S@�ks�J�n�N���a�+{e+�PN6�'�B�7��l����X4���G#r�ʊ6)�6���Bb�֞�D�>�5�����Mރ3�rC�?"I���@��vx�s���'(�?6��2��v�Uy1'�'�)�h�� ���|S+�&��T�O1QUȑ�@}��d��ý���5�$q*-��Hxbo�¢p�$��%$���#Th���U
	�+\�GTb[�quol��5�?�B�R��B%�ؓ846jc��V�����Un)�Ȭ��`�+�j,���,_����}��ғ�������������_���ޚ�q�$�'��6�mf�O�~��V����8Y���"��+���k�n	�)V�Q_�7�	+\��ݵ� !\����19�����bvv��w@�2�ؐ(���̧`ʀ�H�����롂�~�M��ϋZ��B	�HT����ɏ���Od��9!�~j����`�v�n*?Z"��R/^Q�H��o#�v���ݤ"�tV��_˶$� ����|G7�@��	�l�F�1�^*@�7�_ڊ�t�(��s�M�䳯��p�ȍϯyؘ�����kD�X����q�  �ӻ~8M���C,m���q~,���2�u0���5?�P(*����%t���ށ��ߦٚ�3�L�]v�!My�?�X�2/Ҡ�*�v�E���Z-8��J��@I�q�� K9dF� Pa'k{-Qkvy��_���v��O�p��܈Ǎ����$i��
 \��j�� q�	)8f��V�зC�]�0h��iv\t��"����bK������cO���!��fڽw�����j��;A*��׎���Y�ѯ�pX9H�m�FSIG�ɂnMR6)��q ��>�!M�%tf�ud�$�mOl�����ӅZ�*�>F^���e�L�Y��`QL�%���2�(�S*Q�iq>�+��ד�$�6pLm� �ߢ�����8��O��_�v�����&�qz�#�!���7�ʅ��,��Z�3X��ENq�Z��SG� >D�⤆"���ddqG�)�[��d�3��!�0~V\0���b�Du4��tp�0��2�����6���]��g'h��ZW/���kbT!z�j�p�g��&h��:�Hj�f�	�\�܂���§G)g�O+r����#�L/�K�%���ʝ��H��xI� jR�o�P��S!f&DI�A���1������xa�A�Q$V�f����C��i���?c����I��?��)�|���	���%�Q@�R��v1�����zɮ���oh��n,<����q�/����S�)JDg�R�91�E	A���%��`�:Ažx95fϋ�σw��%��
ޔ�-�c\�El���C����u|�,_�K���������,(���Z��d��HӺ��5�!� !_.=�xІ��
�է�n�B-�9������*���^�>1�7a�:Q�������Ue���L��D��=����P����l��	���M��nu;�.Ք�ۉF��Q_G��b+*Q�7�m{��!�>�_�D�^T�)�91�&,��u�,p�˩lp��f�	�=�iA3�L�z�Z�x=F��"y%��:�6s��b����؁�DiÁ��:�+����� A�Y�ȡ��S���m*�.b<�D���������}��x��\7�7�G�YHӪ޲��o�Q.���"K�zql�x>��W�lF��}��(��,�:��$�4�����/�qoŜ��*�1�q)9k�
"�+�H.��D�����*ڏ� ��f	���C	��	�:�j���%�D�8aI��w�a~�\�}�I0<؛Pp<�P���rx�1}�;ϴ7��Vx�T�z�ij�4��1� )ʳܚ�'��8�\�(�����Y'ml���]�p�e��������	�Z�|6��l�oߧ!��H�_�D2r���jt퓡�����m�D`H)o5+9�Q��K	k��aӉ��VHMe��k����uQU1�Ek���v��P�;1t̅�n�r��U,zZ6zaЌ�6�� ]�WW5�B.WS��r����}2YV,6�4A�f��J��-�	/u��
ۊ�<SNs^UY�e��SRS�r|[��t��_7ý<ZF"��t����p���b��Ӽ<�#bd�vg�2�Ÿ~����D!�3HŶٛj+�m� g~�>µ+�h�m�����*,�& �`�Մ�yڿƪm���i~��}�;��
�v�5]��Q@����
7�Ntv�#�V3Zj̓FG�G�FG�z�'C \���oX�iz�^Z��3�l��>w��y]�d�Zh�je�CV�����?�,ʅ� @�_��6:���˙`��	����.�Rv$�4�]���[5*lE!qe�  9�Ԁ]�ӏZ���B��&{lJOK0���ب�?��;��T���LJ>F<APJ�u��/�<ű��0mP�p��2� {��#�&���7c�e�q'�8Z$
k�8;�M�_:k�n<��"�u@C�-YS�	��u�T�S'�o���>!�3 ��+k��{��ג9u��SX%��Uo߸
�:0��"\j�����g/@SA2Z�o��q=��EB��V2�[�Ӡ:�m�-��J�×�}*�#e����p�����$�ـG�
�w��r���`xl]V*�Y�~R��������q�-�#�3	v�p)N�����!�
VH���4�	J;�@�Cc&�V��O[b�f�V��D�c���c�
���TBp���d�������S�
uV����^@�/���ں N��&�@��̆{���Ԥ���D�[ar�x����r��^��S�H�զUY�����<!�9�k=�������܀y�l�p�D���7�p�9�I��z����x�8�Km�����kh]_��Zb����_��0��Q�Ĭ����D�:�/T��ցK��}	Pͼ3�B@�J����-�2�
��{�^�TA�#$0���>AZV-�~s)��c�D{=��0�� �|��M��\����=ۃ�b�?ft�Õ{˦�p@��P��8},�Z���y��ԅ�*���h���]��������H7X�$��K޹j�U�n����:�lF�+"�ʋJR��!
��|�l|\����
Z������uuIo�}��C��g&)5�Ef?�!��S�w���%�U��d�Gz>�N6���\�	�vl�#�˓/��uS�!!vec��G�jj]x��ʐ2�l�� ��"V�8Ln�|����bK~=٫�#D S���3���Q+�"/Z�Ip������!�ۢ� ����/�
t1뛭W�D�5S����qJ(r��'�Gp�6�N~��@��Bf��,�Ϗ��G��گ�� iZ	��;�*Z7Rd���V
b���hnd�~��@�� 沀�V�k��?��_@	�
�E;�e���D-"Rc�e��$���v;�)G��\_���'T	���擻��g��Y�&'�e����ɥ��[�{R��+Ȱˎ/v�W�8�����]|�3b�>,M����v/*�t���v�N ��X�� CwT���{���mc���)��h��Y������7ڽ,]@���)���*J\����9�t�: �Xʘ�2F.��^����uQ�=���		>gM��";��lq�t��Ԉ=J|��=�����`C�����E���u1�4(ԥ�x�5�j�~n�afЏ7�P� ��v�:#���'�!r�\�bu#%��4@i�GF|�g.�W���p��Jv3b���Dۑ'�'��zm;P��c� m��l���h_Y]�9*vS���(G��,M�������J8.��_K1�S;ܢFX�����D�@$e���%e���w��!B�`Fg׫�� �rruQo�~w���Ǯ�$*����-��< GH��L�8�)5�'�AԬ_7�ٯ3j�/�NW�:"�8�8۬A�(�s4�zc<�G$�=�&��ȿ��GER�.���Z���	���gyK�Y��;ͻ�
�3>�Յ��Y�7�� p���r�Ef��m@�[yT"q"����&W��?�d�Ɔ���I�.��pi2O��?b�s#�_�HO�җ��K�Ժ���)��Lҍ{���ro��J���VG�tW�*E�������A���|����]���#-���f�����v{�9�Ja=o���, L�$輲�|M�s�����2�Z�n9�ͨ����(���̹����l��ŢO�J?�l��`(�E�V�C��c (�M�w�&�	q`�1�ل��fe�xs6�3k�곂�^G���I�^:�?0�f�w�.2n,i0�z�k/[3�ҮG+�T�oE"j�_�>"�t����|!��ݮ@�I��Y��U��!���n��j��jV/����
s�4A	Ip���3��C����b�[x.�c�ScA��ID���e���N�'�q�t/ņ!X;�QMk��l��w��U��&�=���Z�����H
�ɲ�=���\ώ(���Y��!u�d|�E�ͷ :�Z����������=��V��;�~-\�Z�q�P�7�Ύ�T������˭�O�n��$��+�?褘K�|�'\�4#&��LLN'�YY�}_:k���%��P^�~�/|��;��p��~�M1ƪ�H~�N�dRhn�-U�]]t ��^�f��ͲU�1�"���0�i�&�	���
�Д5����͚6$l��q�����^LP� �<W͗�U�q�8��R|�1�A]&�Z�2�_�#��l��ǒ�t�Ĩh����g��������򘢽�+�%[�A�C�Y���Z}�fǛF�1;��)�EŲ���L�Њ̜�P$����0���_~��\��c�^�Y��q��K�����$�ٷ���a�rH9�7,�������W���b�8!�m���>���˅�E��֕�j���,��6��d�<���b�G��~V�K��(lSr$>����$� Z�ů��B���yD�J&AE�Wz8�[�lk>e��RG��O��u�:#Q���/OY/�KCm�=k�'�,a.�T���F��7���!7��� �Wf�H�
͊W%�q]�OU���+<M��0`{,�B>?"�����:���)'D+H�`�Z��54�:iIs����� t���E!��J3A�\�g���M��:ҩ�f�pBm��!J7\��m#�����.a����'5��6�����4��G�eo{Kݼ�'�Q,̮���rY�"�E��[
�gL(ܙ��9!�8_<�1���<nq�a�����$Q�"�WC��¿����.2�)>�}�na�{���Ryk:����392TҼ=ZJ�
��?��T1����sG�@00xU*(��S����T9�}�4����ab}uG}@�o�}^_n
��;G%���`�E�	r�0E1y(7�s׺fؾ���ՓI"�k��Y���:��������?�O���k��
��I�`�j�ǻ��+�z�姝rx=[]�9H�n�6�}��kd[�n�(|L_�}�JI��L�l ������P��| ��y`P������$jt6�e!�ۻ*V�j�N�݈g��]���l��n%���u%��d�؋�T�`ˀCt�8k��4������	�S�$ �ܒ�����$��)��`�r>���/�3�֦8,�J��Alm=�Iw�����H�o0�������7��Y� �'2=��f1�~��M����ɣgH���/CʁAb���VdJ�
�y�}�s$����� v��k�G2b���߇G�:��"S;���W�Mo5�j(���v "Qub��z��5�G���������Z�4��@q�s�"��N�ş�9Wý����T�Z�W���>�U����'��14��k[k�@Yf� tp�s	�@��n��J�\�x��9e��Q�^T]�VJUwG`x�BbL��M���@��D��%[<�	��Y�B=�wQ:g����[(�����x�o�V+%���	h��*Õ)���ٟ]�aI�rxY�Y�X�}��������j�uYJ���`��#�rVmn�
�ߠ7Dҋ��}�$��d�B���z�yH�ә�fLP��\mJ��Qʳs����iB.�R1!��;Q-@F�;��� ��^�-�|&�Ϗ�dC�����U.���>=+D� �]o��!3���&c�>J��� Jf���5m���6���� r	B�o�6D�S��nK�ųa^\����̋���Z�գ��]��s8�](R]�`8�~_A�mY�S^�)�.�[���z\ֶ܆��s�p��[;����I>vy�񣠤f���ɷƉ�# ~ɫ�8\�pK�����d��S(��Pk��Eӧ������{_�s��R���κ�ǤMI4*<���W�B��U�O�@�5��l�噀�Ѩ��J�=����xo=����U����G����Ղ��'*��+��0o����@T��͠��}��\�s�𑨲���zg���tJ��PO�1��3k�uvK�|/A�?d��m�RϾ�Ҹ�:��Z x{�+5�������=z�zj�&�'6�"_BZ���;������0���w�N���A4Eؔ���z_�nR�1UL�g_ ��`���6��;~�
�7��Uڔ�#=�XN
*0��H�1|���z̅�,ٟ�z��ʋ=%{���� �B�����'UY���<[`�p<�uҮ�$��=�j�0�N��t��1eg�U��fN#z� �����M������{Y±�������[�z���+�t���;"x�-!�|>C�;G�h��(,k�'�����o���K��M��T9�r<2��Oȱ�WR���4�;��6MP����@i32��)�ة�� �,?��nsއ��QEf#����a�3�@��D���L�!ą1�rs�	���`�^ȟG�T���̺�aw6w�zO\���v��| �*3y�up�`2ٟ�8�ͳ=G��:�D�\f�-hi�(�4�2eU(��F�t:�m�.a1s�I��f!%VH��pe�@iK/�j.���D`%X����n���ґG޿�H�� W0��i�
��od�����
�����a��e�b���D��)}�ΰ�V�݈�jˏ'�A�u�a*@,PըFIy7��P����7E/tA� �sE��K{��?��]�`_���p��j��be(�<�.��uЀ�e	*Q���T�R�!�&-�f�*���5���`�B�Ϲ^o���ݩ醥u3|��V����	&�#-Q��>��-���HB+ס�� �0	v�p6�YH��L2���H:�Б�1H�V��!o����3w_�n	Ԥ�7��{���k�*�B�T�vd�y�Ξ\je_�����Ԃ�D���T�����c�%���eۛw������G�S����\�Vw*t��v�����@Q!|+�jU�~�?_(#m��a��n)(��ƒ(�É��>1�k���ٛ����%���Ў��� �`մ�����Vل��Z�� �I��M�Ll��X�gM��e|]��MC:�-0N��L��+Xi�gՌO����"��^��K�v
k1{a���0޿��;h\�P�5+�ie5P������Lʝ���x~�i}]� K.Y՜�j�U>yuj����8�Ȇ?��B3VS�6���$�k��y�J���"y+��}Y��'4[*�zy�;hQԯ��5��L�=Q߲�y�NR�hf�t�8G��D�V�q� \���_��՘q/~V9q۔.'L�7̥����&-�{4�=�����
��H�
�Y�mK�"�~��6]״m�LW;�8s������3�B�s�H�o�gq�L:��Zp���0��5+BX��i�M�!��e��H__�\��[�fI�%�.ɐ������������I}A��[3��W(̂/I	$��@r��H�g��w�`Rƌ`t���@�D��2�t8���?z��ӿCߘ�q8��۠40��Ɠ�)������]\�t+�I��)9>{!���(!Y~Uo�d  O:�?��9~y��T���1B�Խ���)r0f������粵�jg��K�����on�%Z�����!C�p��(��U��A�M�GV����<�۹�ԟ�)I��S�K?7�
�_x>��(�L�ˬ1� 䑬\�MD?���Kk�2#�y�/�A4�e����`x(�`fXw;^t��3�hDh�����"O z��Ű�Ȱy�%�ԓ��l��SKq8�p��șv��4�`�U�ނw
�L�� �e� 7�TsO�� ��{�G��w�%^�K[7�~����2��� �����]7�����ɢ��05<ݦU��`m� I�\X��{�C#}�uo���0L�ĥ��p��]*E���'�<Q����)WnXk�m�ⱡ:��!�b�G�j�C_�cNZ�+�0�[�R��̈�ՙ`�	��f�I��y�L�R��v�7��C�V��
xm7:[Հ<"��}�m���eߑl�����K����6p4��k/��qX]AQ:]�:�:�m/]���u9�:��Fź8���_�=���3�#�Uؾ��
~D\T-��-m#cOϖ�ǉLe٧�lYӗ�Y�3��n������	�0��H1/��P�y��4J����)��q ���k;+����Ѱs]1��iY���H?�WM��uצ{�cr'����
_�hm>�sz��v�������l`n8Qr���U< 
,�Fv,m1��e #Q��&�����nM8"q�񯖭�r�U��D ��f}�'�����֕�S�I5pʴ�DEZ���-���3��~6��ȔC�J��;�iEt�a�P</��L�y���T��w�7�e{�+�龚%5P�m�U�Q��Z��U���5��`�MUqc0�ǾP�
�q��<r�ڂ�o��q��~���d���Q3F{�j7���gW�1U��p����� ,cQ����Q;�܇I06\^R��k��L�-ƀ	��7i{��g�Z��� m�f>��<&a�7 :��#�h֖A�Kw6���=�\���ɚ��<��n�����m���[t�M{K�Mb�ޚ[�黙y �/�d,�D�@ȭ�b�_&�ʭ�2�P�	�ud�}�=^�����n[Y�A�L�ޮԚ�8�/�	��'<��S�C�ld5�[4��|�t�!��S sm��v�?����f�8�-��(;�T������"E���i���`w��,�j�)Sx>r�v>��d�n��b:z̸+�L����_~�q)0�z��O��p��w��wb����[-	3$9@��_ͥ��#�ǯ��6�d�����+�m_��##EA�����A�4�4�~T2�5�d\�y%O�$�3��"�1I/��G�I�6"+70�k�@�	�C��^ a�#ev��-8�'�ӹ�?-P���#�x7�-�eakݕD*U�Y�@��:�t->80��+W;ʅ�S��!'৘S����#�����o\H�g�m@j\G'J�[mwʇfW�o!��V�Z���O
�)R?���T2i����p�Xh���Z���ـc�?X�o�ʟ';�v�^��)ܠu�,�aaj6SL��WE2��1LS���FH�B&�����^��g�i"rC�v*7��ߕ�/j�-��׍�LpEާK�̤�E��YMMb�JDu�|ofꋢV1�y���0
NÌ��%�A��xͤ�d��I����( �
����v6�JB��%&hU�%��Pzs�|uO��H����S-�ZQ	&P�����i(��*�Db'E`8g�yf�,��u�uc߅�g�^|��H��\[�gX�h�/�_;�6��؞����-L��t;�eS�0���e���?�� %q�JV��� 5�Q�:�"d�C:���T�"���J^=W�;��ob�O��y�	�Kd�-"��i_=���z]yN�X�c��F%jm��:�F�>�?�HݞN�RL�W͍�.�{k>})����.�h���ō˧�}��f�o<c޸�d��f,Ҙ�y�Ɋg/l��_�u`@�e�����g˟����&�
�:ö
�7=S����F����D��ݸ	ϟEEgh����U��`"�0�(pz�y�ɥU���!���l��kN'��Bk�����{���2^iCB�L�JB�i$�`3�io�#/��AI}�?X��K�ٯ {W0%5�r�]Q�'Z���/� ��r:X�����5�B������FFŰq�^9�mf���f����{�o�Qm�E����/����	n�e��(�e^z���^���7W��Lr$�u�a�iH �
!aHR1���?�*����~�1 t4T'
,8Nc�]�c17Mc<�8P-�~����
��B]=;��&�  ����oc�MP��;���璃��7�������Yi%z��E���vHa4D��#�֊Jթ���l�7�q�J���Pd�.�%,�G1"�x�>(Q"GŬ*���X�[^O)7�]�p!�*	Q�2j�vو�~2�
*�z��.<�~j�.���.�sX�1�����%W�.;J��@"����B-g��ja9���A��ca��^�v��#[$��i�"5�,�|�|(z��D��_��u�7���(��G4ѧ���
���^���j,w�I��as����\c9�^ı;�3�g�ê<�`(/������8��~V��_9������)GڇؘI3��~�����M`��P��C"�(�9i�~�v<��'�F�!�V��Zp'�n�ͼ�����^t��c��S��p�.ڥ���6Dd����Dߗ<�*�̦&Ɛ�@(O����+}�aM��@c'n6F�,e��b�_�V�9j�wnl=_1#sBaMN>ʪ�|ƫ��|�vT�PE}t�V�h*���;{i�ͬ �T�lBȴë;�٠�vPP�R�@5�esjF�nJ]���a>"�;{�m9��BX��E�m�y����i���C���3��t?(���#6���%Q�?T�e�D�AUm0&fO�!3A2�1QUR�xņP�Ib�[]wV`�}DGD�m�je�&[�*�@��&)\�V��?�{�R�8J'��Ӵ�t�(r8B	C�4a�H�?F����q,z��1�.���k�TO愂!�ӽ� q.��d��o����ˣ�ռ2E�FT1�ݿ�_,XDO3	�J*��v6PO� 5fT{�C�nCR�7k�Lj]4Ia"�L���s��e��b�W�����c�Ș�������\ᥫ�r�1&�b̶���k�x�z{�h4�b2:9��Fä�:"^2����9��w�(DE������%jf��K��|�R � >�pb�ohK���SI�v�^�>6\��u�D��\�@.�ϫ2�ih�TYH�!������%�>�b�˹�Ɓqܔ�Gl%M�r�-��vPl��;�:թ�".0u�=}(��r��J^�~��W g�-��n��z� ���0m����5W��X��dZm_J��z�%Eb�ы'��8'�w�Rk�l�)�(��Sg)@�~+U)N�_��J�b�Q��()�� %���q�1}�>��I��Ty`��*��?ɁPq��{�e�G�XI���	Y�G\p(Ҭ֍@Ű�M�6,�0�^
p�����j!}A��岫�&pu�����I�6)�ݺ)
+��ӽ���	�&��B�gl�=�>��ɰ/?4\ܥgz�7
�n9���ߑ�G�>q���*q\,�a�]��\5�'���g��a#�@:�� ׊�Wf.����C���'��窺�{�q�K�*�V�����L�t�̐O���s_��.����@r2�m����T_�����@K��c�u�%ݧ�	�![���
�I�4��η����=�oՔ�2�[��˖�Z�@� T�J�������b�}U�^5�,T'�����`����P�}�����4Ҥ<��O-Q8����I�?"��}���Զ�%Z��(ڡ�=�a������G�HgP�T�|X���d6&[}���d�k�=���f�	1�p��N����TOG~��	�
��$z%�
���͍
4���o��g�$�U�K�/�e�4X����:�6#��K�2��;"�����Ni���N�*m���p�l|�Ƶ%����=V��Ie�4yǬ�"��(�X�+2<��i6�OmR�(��n��Z���n���o�#�Q0� �-�]��@փ�6n�c�/9_�%��h}.<�$S��}���n�u�+�>a�7I\�=F����5�xٝ������a��Mܓm��í��]�0��)9ϣ�QB ���(��=S�{�5$��t|H`�t���-3~&���6�i	;�>L6M7��()x�hn��>s��$��K8v�~BnVG��nDf� ��3�Ы��b�\^K
7ʷ�^L��:��5��*q����~���W>]PD0����i�� 8i�]!��Y���Fw������Ug�o��{M.��1��oO�c-��#Pf����&ޱr��"s�Ǧ�;3�w��F�,�<R�pȧ��i��5˾�
���j��k�9��e[#����ڔ��s����Y�eE��%���EJ��,�$�:�	?P����ɬ@))�~!��Ľp=��xAm��z���ku�)����G�O* �8 s5 Bp�P�s5�̗kx6<�9��I��������x���9�*���Ѣ�a��8��[V�B��2��A�#H�T$K�GG��K�8Y���Z�n��m�!r��Mx� ��S�Ql���X�#�N�7����.�e�T�3�᪽4C�Ş�[=$ӎ��MG��*��`�d�}�OW��m�@R�
�|�6���~�Ϲ�g� \�G��������"K�'��=juD� od���*�eL�5i�lW����� pf�?��d麼gY�����mo�,��h<��^UVQ3J����1�r�Q{�e�v�����B�'�ݛ�ծVv]1=�ٔU��6K�s�j�!��o� {���"�ޥ���}�fUd��BJ~>C19��Z�~���w��/���,�����@�y�<E��m���8�܇�=f����UU��l��]���驊��;Os5B6C�>;�Dڌg�B���&�#Y0h�Ҁ 1nh��|3�5�n�S$ų�x��id� n9�[|�4��7�8O`��q���ghAa��=�!ùR�����	:o����{'5�L&�c�MP?���Y�&W��d'��7�|�<��g�HqPz��6��B0R��o������B�<�J��W.�aԇh��ު!R���?Н�����_��f}�T`I�Nf r0�L�	����Nk\}��<+�wԪ���HG1
DHTIRj�/�9�54U�kSݲ��`^z��vqtʋU�-B��G�ou}�p(��ֳ`�481֙_�Y#��i���/�E̾�
/B�E�V\�����3]g���v����a.�=#�쌹J}�}�P�j��)��3��z���}$?�3"�p���Am�f8oj�k�u�#�!��F�s^qi���E��fg� �<���k�Pf^��о�^��nU����@�d_C��%k��9/��.UQ�������� �>�2���n���0]����b����1\��e�Gٷ%T9�h����6�LB�W�)k�`M'q���>zX��t���M^G�����a�nh=J5W�O��/�$��`a���IX�A��}���u`p�����'�Qi���xm������dդ�3�}��,�5"b���}�+R1� ���N�&F��9�D�L���L�ې� �'�#S�e�MنNu��p9P�4D�����){�B���_��ybH�~�ř�|�YB)�})��T�م͐���ˀ�~������j��ԅn'=��gcm��>N߷~�]�N�����Ȑ�w��������{���er��OW��mfJu��,��rc��6���o�	nJV���T�f`����Q�SI����jYy�)�I��4�B�i�;�.T]l��jF5
�5����֏������j�g�.9pR��OҴʴjXa�b󯿩��q�ǽ�,���L�L�KUbq�@v��$�֕@c.h_��(�M��w�r�d��a	��̟e<i������j�
�^o (?�P�)T��Cǥ�� �0G�>�SC�c׻�7�dE�f���ik9 ��25���<fD�ͻF��!�'�%c�l4�yӥ��	d��ur8��K.�e
�i�p���3�~/���mG(�C	�>���Ѯ���Ҙu^1�vr�H�O�y@:�
/�e O[hO�P��*C.5��'২+�Vf�ݗ7���C8y�^~rg������Ύ����9�����E��ܿn ?�`�xR�%������@lSKq���!�L���/_WҖ�w��	D��/�L�яpH������q2Ҟ�3`���T������ß�n�,�˞dL�QOT���/��v�,�z�ۧ�e��1P)J-,�럂2����!�Hԫ�^/W2���޺���
�"���\0Y	qZ9:s_غ���!d	�JF`�@����p���Oc�ǣ��7+���3x��h9� RĻ2�͜�a2��0{��e��eUa=|���O�t���{6��9?BCIClx�-�� V�8^��IW�y4l)�w�~"�G�9�B}��N���F��J-��� Z�V�w�pU9|I�bQ�����H�Ȃ��������	ڐ����b*/4'f�ٞ%g��$�\�0���$J*�����rs�?�!��	f����V:6�n:YTm���ށ�W+�i�u���'<0����,�*�hV&1�L"b�gl�D'Z�����q��$��#xߢ���qI�w�$]�Oo2��Gj	�߇��f�ޤ,:���'�_3�ց G�
zc���� �n���*�@$�}'�G�5:��l�@��;m8nȎKM��Z6.:���(Ұ�3��)O��}H�bl��(��h)�)��������B����cTR2�j6��w�?q%�#A�IN
��O�GV�H���ׄnX��$�R UsGU��*���Z��� ��[ɉx��P���,|�D���3��-מ\�9�ܹ/�D:�m��a�1!�Ô邘���%F,$�����E>���v���Td_�@���q_,�m��)��Z�ӎ?~�%��S9�����bv�]��K�9����ӓ���+�&���`��T�I�f�)���0f'�OA��C�����$�9t:l���M���L1�4���7ŕyi��qr?b&�~���Ì�^�L�:+Q��2���7��`}�H%��!���cf��L���"w�d�2|�aB��UN]Š��\�H�v2�g����]4�e���P)�nFJ���}\����p�Ty-I�E��|��K6{�馧Md����N���#�������AZ���a{�R������x������t�?�u%g�	*�\��$��RW!�W�"�T�d��[�fo��8�5 �v��R�n�I}Y�#���t����,[W�ܙ��wCUt����靚���Nq���I��Z{��W�V�J�y�q�Q�`Z��[`�~��P���nK;��z]tm�-0"���V��cƍ�ir�f�U�-Z��iZ��ZC +	�"�_�X�/<�$BM'�� S����^̌o�}�C�X�O��
����j�S�Pߨ��&�bϣ�����Խ�H���Q ���H[�A0O�v����ҙ �_��(9|⸿��D�"M#�3{�&֧��~I�?��7	��7Yh��eG+B���'�գ�X�Ec8��js��{���<��g��ӚLN��΄�'��Ʉ>_�C�$�Oco������whk�S����u�V��;�o\Y��d��3I�[�d1�3�h��6���>'4��|E��n�����0$�k�,�	'�����gO�9�t1�_��K8;��P��J�b��3�F w�ƌ=?r:�b gk/��_�G�f�c#w7{g�6x�~?�f���c��R���ԧ<���~p�]�5!S�]�l��0+
�rB�ϫ��hTg�NΪi�l,�Cy	뽗(����hE�Y�ݾ�������A�`���J�;D�.���E��r��7��𖮙l�׬6�L]P��R�M���`�\��G��1Yj�2тcB!���b����-O���������K��1�����r�n�rGv��|ղ�o\�^���~�x�3N��֔X��2D'��	@O���~�G�`�H�)�M5���N��?X �5���R��&֦�=L�N;
Y���K���!��߶dnP���	� �MU�Vh �A�;¶ �ړ�y�$P�l��k���m�k���	�l�U؞�^�_U���6J��T�C�~	h.i&����	�E�IC1.ޯ;�ύ��ɊP-����[K>J��?�D�p�W�1�rҼ&V �@�˾����T��2�jSR��N�����E���?�'�Z���8.1�4��k�r`|��V���*������f�̗�$f������MmVi*%�9N+���Z+t��p�|:2����\��a����ZY���AE6�=GG��A�7>��M8ЧrI�䦴*c�r��@�W�;�@w|}��	c�UPي�)DKSV���a,t�ωN�*����/���fל���hr���Ф�t��:~�q"jٳ	�:=��.��S�}�?���-�4����)�Q���sV�5���}׈��:��NRNr��G�E�%�-,�_[�x���MV��(0���Wkmgf��7
W�2�#�^񑵏:���c,_�uL�#L\��封��.%�:����44��"�(��7QT�N��&��V|�ӷ
��f�D��{�8�5�����v�U)؁�2Bu����}�眃�>
a@���S5tO��֜s�
Gq��N�k.��Ž�k��{��e�a*����(*N��ʮU��v��z�yoZ��
g@3JA�S�J7%��⦔�܀�������"b/��2���/NX3��2����D�6�fI[�����]��ڇ�
��/BF2d�M���b-\/�@��U�6>e�j@�4}5h&�,����l�&TU֦ͩdd�0A�k����^m3̚IP�~�\}�+�#L����v��o�W���X��#fĮ3�?m,�t=�x�]�D��Y�R�Y�=/����>eK,�nI,�b@�ڄ~�>Y�k���Xb�*���&�̂_��%:^:����H���ዳ��g��j�
�+��{������uR���؁�$s���lz��\�l���X��i�~�X��T4�N��V�snS���iK�oT�;���hg/CN���O�D���M�a?��Ԇ?��ԏ?��H�J�(j�˂ON<-w��ޭ-�Ғ[�ȟx��^�>��* }Ň6,xRI	,�ڜ��a�u�bčȎ�D�~�L=S�wV+��w�����$�1K����И���.?�a޺��BT�Ҧ��v� �=`�V�K>�|���S� �!(����'۶L��E�2���qw����k�}j=�r�F��ƍr�r+d��U%X�5�C�;&��M�ʚ�3a�#{�b�
a�P�5Շ���5���'|j��_��bj����ڂ��Ʉ�5,�p�c��=�Utˎ���ă`�>�2����!BV��:��얺�H*��?&����ڙ�o�/�������,w�k�`v��#]x���&/̨l���t�r�;" ����%-Un�b:�u$`R�Қ��Y}~�F�k�<�+�/"��� IT5��U�XZ��v���Wo���B
����>E�, �����l̞G�O]]�	�F��{�V�o����u(��e��	\i��	�H� $�O�D!O.��?���_�w���4޾�Y��˪��0$/T��εCP�{m�
{h~��2��v��;��w�G�@�f�{6�g�{j�F��b����?��l��h��?��	�$K^�����g57R�Ez��8OH��[�"�ݜ�[�������_���p�����{m��(�%��W��t-�[�ÑE�<�p}-��+���]$B��m~hd��
I��'9Ў��w�{��{1:ӓ�O��D�#&W-�%3G�� U��}�����Ɯt��6m�.��7��~�K�x�.BAMk���m��MA��&蕠�ⓐ�Rx���,	i4���O�i�hs���	hR��%�N�ג$��]-^4 �~��%9�7� QO-��M�^t?Z��|�l��G��1�]�Ȱ��N�Q����$S�!�n�k/�@0H�f_�Q����%k{���+�T����p�Jm\��9�K��%,ť�~�4�ȉ�4�}In!�R���ĝ޵8LSt�����	l��gc�%c%9�jg���������zD�xs4|��G�=Σ8������/0�Ot�f}'�S��3�K�@��͢ܭ���?��^&"���:]��F(8���v��Z̞ood@R묷s���8�j2��Fxc>���`�8a�p��(s� �o�d�r�@��3�<
���uc����b�䗝!wak�;��G?z�,ߪ)hr 3�����udW�X�|��9�>���9櫍�\'�Q1�%:�VK�R��+m�� �hoυ{f_<����a5u~�_�U2���L����5����6�1K���z��{�Q��X5�,8�|�",M!�T�:���Y��4�h ,c�r��%��w���x� �l;�b��w���8�:��'����D	��D��m��3z�]�t����b�3�p�W2��?�A�9��Ȉ?2D�$��d�L�-X�m�N����"W�i�<�9Ͳ���F>��[\o��d4�]Z4�~��P�v�`y���J�5~��~����W@�s���{���yz� ;ړ�wD�q%�٥[]�~�� �FH���T�T�:l�n׻�>�G`>\�Q�%����8KB�,��b	2����(�e��=6%6�"U��8xW\�ù��p[c��I�b�X��l���.,���Ih���TvR���� U���d�
�j�W�M�d?+Tb�u���r��L��
S���URS�.T��HB��>:�C�9�і�`���,�0dcn��Pv��p��w�R����F��$e?Q���+�N�@�����N(����KQ�� rqY�U���\qWv��CO��cԅy��B(7Qg,�]Z�Uw����`�J��I�G���+�\�U�,TMq"*k ��sȱ-%���(e��~�-ߵq<Vۨ|�xʥ�L�|-_f���J�s����Z�S���7C��ö�3
2X'G�蒽�=���3�x��6�"���Z ��	�UdF���"�{�*��ʱ^��Y_&M-i�K{��ﴁ>�	`���S�l����d���5�<����6���^+�k�+[@�a������Lvu�G��@\v�j��m�B+C�CDJ� W�z궩Q�kh6o8���vb(c�pI�G��Ǣ�?!�}ʹ1�'����c<�?pW����`'%D*N��Y!|���zZ��5TF��@���,��8h(�~����&�����i���16qc�U�_�XI.��BZ)�R��²'3H��xkH�PxX�H,��{����c�⨤������T��h[\l��\^s����q��a7���(�jz��T�I���ju� �R(���}M|�:Y�N���h��c���v<�g �F��_?����h=�mT�^�h�X�-�����D��rQF�m��'�\A��BR<?�X�:�oO֯1n��q�]��1��2s:�,v*);�b�T����_Э�L�MTJP_^�܇#�'!`������dለ�^G�pC.�P�P��P�y殸HNU@��ԃ9ڰ��A��գ| ˩����Xrko�"��tT�_4�ĝ�� ��M>�\���T�vް��<���(�5{��2Y��$�n�����Q��e���"b����}��cǻ���K�+�E�� ���s��|�~�I�ɂ!��lT�kS�{ryz�T�3cvR�è�D���v0��\E�К�5d�5S� )�}�+�%w�[v�����W����m;�3=
�����n��v�:�7��KJ3�����������F\�yb'��<��w?�Tj����:9����-����+�&�CT�M�>Hq2@/��?eP+�G���W'Y#6&Đ�TT�8�:WsNH�d��{��]��gU_.��uHE�,����c==w�O!Ԇ�������s�8I4��/���B���R�\L�t�e���t�ð�k����z�W�IM$�d/+h��r����2�i�ʠ�^~}��E YKQ-ON��򒚢���(�O.��\��a$��_�	6pGa�X�)�ט����k#�(%D�Χp`�#�t���F�k؊�U�o7�v��t��@��s^Ŷ��-�[;��^���B��`��s���Ϝh�&x�
������~l���S�H����@[���r�����W2��N1yj���T����@w��x�|����P"���u���f��$��[-�#��6� ���x�@��ez)yPu7��������/b=g8�q�Kfe8�P�6=.�4�5@�nV��]�+��v.�
��m7-���L�14!e��f�քE�(���XZM:�}�O���QY��Nנ:����x����[�:��es�"�1x�L��lf����yH��~7���1��i��W�~H�r{�׆�?���'�,�[u��.���5$Hv%6�7����n~�G�AѴ��F]���	t���{(l乳6�s���gt�0P��eQ���	^��0���؏Y��b� ���G�0���"��O�ObT����{�r�WK֏L9��s��9�U�.=�,����c�1�mӍJ��� �S��E�i����Es�����(z�u*B{�N 2��b��p~7�/���A��J��ךm7Gł��C/d�b\Q6�R"�d)o�4���M��N��twU���o�?ʰX�σ`t��1g���:��Pr}�t[�.�1�W�x�W�V/1׷���O�R?�Gڻ��y>�Y۠94�?�b�tTӬ�07`-J�q�R�)���Xf��b�� �������z��Y9�gHQD�X�K���n'�l�pr>���0�Ӯ'~N�P��/�-�����\fQs����Ŧ�vK0p�{�&(����p�@>}����D��#{'����6w���!у�m���XR�a}|ߖ���oܭӑ��0	Zz�^������Q�<��ɏ.�PV�d_�^&<�F��-����`ұ�b�����h`H`Mȶ�L���K9��tϞf�ՒyQ�Uɉ��ek؂�Y�OwJ�3r���0�*�����/�"�ӤOY��2uL�BH�Ȍy�pw��]C��X�f��S��]��dNu
b9Z�֟[h��V��$l�Ka�S�����^�wq�#�ÒS/?+�W� V�t�����{��Y��[��>�:����`qsJ���Eh�ۦ[XԔ,���lx��26�Ogmt��$L �����QZ]�/�f-��>Qb��-��9"<�n���� 9�WjD�i�#��6���+��K��?ޟaԆ���u�y?G���Ѓ��f{�35<�^��ɐ#�;V��&+M9x��|1v|���sZ��z�R�x2/o������Y���=�[����[��8�@����=5��%�NG�����c���U�$�Ѡ~����,F9 R�K�,_Zk5z곝�i�JM�+�L�r�U����=n�ޮ�w�m�*.�i���b ��X*��O!g�n#$Ho�	�'�?e�қ6D����6d����3��N�7��������F҆]�W�fA�N��N�Nū�h�2�z
�ω/)�?��HTP�$L��k+W�D���r:OL��k�K�q�1k�>p�uŹ=�>�U^�oX^� �S_#=�0��F�t$�-���p@�^2@o�;~c�æ{U���Ů�#���x��%�^7�9v�x:��[�K�1֟3�g��S=؝oV��Y�&���Nsz�8 �,��5�w���Q����l�"��¤���0�����
B�f�D<(<�o"Qd���,��a"��im��\vŎ��Y�~��$f�����K�_�bo�3�4,��ܕ�e�yHC�$\�̃N�,Tp��/�T�'l�˓`����|���H����\4�����R�@�4(S\�ؾ���!ɔ�gí����
�n[�r��i�� �{�M(yİ��W,;�J����Wqǔ\a�d+���4إx�Ujܻ�T�����M�x^���#:@5>���Q�Rf˽�Du���k��n��;���e<�ۗ�r�' �RWlp��m_�3FH�vO#u[��Fy�y��CM�����l�#��Z�3(��R����~5�J m_�}���L,�ͪ�Ħ�A�Ā�o���L3�	7)z`L��j|Ż�칤YEW�
Th0��Dw�p���w�{0)�̓։6X�jF�4�R�H���_�b���Q"� ��U�@��������!o�6h�r]�롆��:���ʟ��6ԭ�C�<,�j��s7��xqH^�?>�\�b% ��(�z�%���?�l�P�ܖ\�Y����L�3�W������Y�]���!���s��L���.E�?�邭@'c�����T�΁w�||�lvIո�l�jA@�Qv�򍭫3<4�)�0"���q����[����QB�l���X��$��uj3�ț�O�_�f�~�s�lr�J*�B|�O�n��'������d���ܟϰ��U�82z5��J_f^e�+-o��-�#�>4����K�L�&zAr�6B:��x�Ӧ!��"p�X3��lo��*mW
��<���!a���5�Qe`�N��x��?#�һ.̯��g5.'%�~Ӹr��@���XeV�GU$��K��p�0��=%���#�#��<H	(?`��6�c���ߏ�����c"���&��ԥ��֕9К@�mR
��������ݖ�5է�*c�|y���� R%m�s6kS�c�;��V�|�/"���	�����d�����V��x3wc��442��α�-�2Ǧ��D��㬄��f�P,��/Г����F�ۍ�Ė!Ρר��9�.b%����#�N*g�q�ÕyS&F��I�R���C�.��0��a�U�:9��l�f-cw�6:��3�����eD�6�s�Q����G\����@����ה�Ny���%N��yP*m��cD�����������R�q}��C�tͰZ����~���C@O�:� 7K�Q�o���h�SR�`�?�T�h/�='f��,�P�Y@�
���TuҀ��x/���Gr���=��P��)���V�`Lmxt���`�l�u������x�)��k������P~��@ѱG8�tju��5_)���%�BH��es��ك�S8�#s�t�@�{�ب�%�n*��19� �ᘢ��bd�DtIm�����D*��y��{L����/ur���W!�]�D3���|h[�K�@�ai�|�Û�܌<B--G�;�)�� �����޼<�Xa���Ew� qw�/��s�ڶ��G�+����KvI�ym=�e���\`��ҫ�Y��0�!!|��"�n}נ��(
(JlX�Ì�*^dx+�΃���|��Rd㹁�S�����:l��B,|���,�DW�Is�+�۴Y��5`9��C�����M�����[��{|ɮGT<��M<�j0��e@��j���(�hޒ]*��eo}|�Ku`���t� \��h�M��T��to�O6�U�$$��<1���j	�0i0�I�F`8�����c�%~ul� �U:�K�A�]_�B�]E��ئy��m�Qo�HKI6R�3�g�?�����0Q)e5�ΣкC��@[FN��H��Ej�\�+Ϛw�i,�2�^m~��#(jsT���#>���w����:!)�I�w�)|ИO_��[+���g�I���rmO����|��U?|�鸏��:� ��j�8d����!�����M�q�N�!�K��j�Wa�7� �gr���UcԁW���4v�&��r�����ho⊩P��7]��'>��ZԒ�Gz����=ľň��~������H=h8��q�H�-��C�^��������$��*pt7^��t��v����4���l�  ^@�!�j��t�'-�r�k�
��a	���2(�
�bm��oeu�g�s����Q���۸���ոQ �W��
��^a�[Y��� �~/��0N�[����m���Š�� ��O�	9�|L����!�a�֥Te-�!�m�A6���q�'�d'����ҿZ���:�.e�x����no�s��\�5߮�3��f����"��d=	�z:�Йg���I6�0�C�Ф�_x��
�7�״`�z��mE-QmoŨ���Q�1�	�c���ډ�����r�:�����>�������Ŵ<����v��nG�]߿I�һb0q�ST�����Z������:-Ԛoh$�hC2��?���_F��y����j��K+�5�	�6���L��fת�fHѲ����]=,���
�9��=O=�H���4̔�s�^���[�f\���甇3�<�m�����̷��7x�Z狓��ɴj�^� E�Eq�4U�����K�e��e@y#����4�+ wM:� %w��ہ�����b�[���_��aV���B���ؒ�؝c��I�C�ަx妆�����x�.�~wNs��G�i����?���'�/ʭߟ�0O}��[ƏE���=�K�^a�x����ms��#�@,�-X��!���/^%���������␌����M��Foĕj)�"j�����@n��gy�}j���l�~w�e=U�ܰ��{��˶!��p�4Lm�U^B��W�.�X5�V'p��=n�f�̰e�� 7�h0��zR��)�p�����tV�˰S�u��(%wwd�CL�IM��@/@~��q�H��)(��L�'I)�C�3A,���Rɧ���*�_&�w&�}5��c��٣n{��)�ج'�^�Be�z��ܐj�7QS���Hn��TO���GB�u%F6b3�e��/�2��{pyS�S�Z�UpՀ~]�@'�z=�-v�^���- D9ch�(("h��B��ɨl��;Q�`f�A�;��v�Of �h��5�.�s��)���j��1��(��L�]L&5�|1=61�]���ZߗN��H��D*�Y�A�������2h�F��z�ybr=�v$c�`\��6�S�DV�L�n���-����G��w�w�r$�M�qRH��b6��>�r[S�B�[Y�����RY�a4�8���ip�Zw�� �:�b�e�����X"��c3f�pS'���CR<w;��;b��;��{�q����m�
���Ch4?"!0��LV��7���}�&L����i2��͸jH������0	GzAU�����Q+�Έ�-4R#����W'9Fo>c���IG�[��O���1���c&]ā�-��*�#����>*�x#k����{�������r�{����F����>"�DHR-��\W`�;�f�����z�}JV
��CL�O-�VO�g�y�2|)(�E��$o
�? �ڤ�#d�si�C�U�]O�Ϛ�h<�T���p� 	��z'Zk�� h�U��^k=C�n��py����<�ƭ�;�f:s��[{�7�;�.�����z&4m����B�U���W�m�Q{�M:9~�,L���#J�%�ܓNDn���?�9���:?����U�)�N��\6%H���h4&�!�|�L8�-��*���q)Y�tes%lۣ�����*qq?h㬐8��<Y�V`�DR��W��P0�gM�� _*�H�	����׫�����H�ن���c�l�5P<��y��{ɔ�ge���U�8�OF֋g{�9�	��P��L7��9E�?|���LZ4�=J���1��m����ß��9J8�a.�tFm0¹���/)�?Q[��ʠ:��V��2Å%���v�wdm�Mݯ�̥�v�4Ns��Ĳ��N�S:��]jw+rn?KŖ�W ��!`1�9��W�F��`OF��b�k��;[�2�7&��`iSku-����1�'[��`�D�ęL:���%<�*��X� �l�c�B�P
;�>-*�����I�����ԥm����.B��l���N�PK>��\�D�P����*k��'��C\��e���a��v�D5ݔ��@�e�g��-k��%�e&�A/�W�)^�6�pثx-+�>浞d�al�j�6���g�����BNT4ʤ��Ξ1���JPE�����N<��i��^�?&�_���{�@*�<N��g�6�~�c�\u�czL�Κ7r������;�%І
b�!YS�
.lė��ҁ*I�~���$�� �.�R$E�.P�HSڡ�=�Le�ܭ��f�٘aU�ŇDڧ�y"I���K$�H��9=��G+Bg����?�YH��5��zq�F��6|b��2����0���5m_�� �+��A��7���^���������?R���i��Bf�%q��hn���`�n/Κ��HWfw�J~ψ�p�m��T�H�t��g�)U��/�߫$
�\�"���PM�(H 15�mK�
%"ua1&P[�!�G�뾓zZtXQ��d��O��5�@��4)yFrSN����.;n�7�Rp��vd�Q���W �5x/�yD�o�9���P�6�1a���$a�A��E�
���VLԎ�(S6��yu�O�T�v������[!�v�oOwdɢw�d<t�R��}W��3�&X�bBv+Y�op��#v�2*�����������{��?����<��b�`��.8L8@ʝ�H%�V,��W]$1tpK���T;F��r���ϳJ�n�k�?�ᓨ��f�KÏz�Y�fP~|Q�.��F׷�������}�E�6O�2��"+���I����d�����Cp����s�'�N���"�+W�A�F��O|ŉ��l���7ۿ�!WI��_=Xj@`��H�q�����yݕ�Y��W���?�y:��>�Vͤ@)WeG@c&kﺭ���)S�ɲ��"�� Q{���8�'�b��#�ry,�f���ߟ��=�6�L�IY���!�o�lS4I�׆x��
7v?�^.��(�t�x��f�=�@(��,3�r��Z9�,�s���\�>�c�xK�Ռ���1[R��2���W��`���`�G���34�&��t¬�}	T���>�TZw���r�<�a�ج�I���D݅��f͉z�C�αI	��'Vx����[�IcKˌ}*�yd4��ɺ$����c��o�(�
� 3yK� �Siz*���?���R+��=�X�����@Zv���BQ�j8�Cڷ���ū�#���*�8$_쪦���LR ����5�h,w�B%�Bvy��0���8`3T�6�_SlYKt!�\J,�ZD�K�G��zM�kX)���.�,hq�N��4�1OC�2����Z91�x_��	���gl�O�B���B�P�S��_�.�ɂ�ь��8���7.Gx���V�)i�Eu��q�	�O�M�:�B�au(�|H��}������?7�L���Z��Ho�6ܚ��<Ύ�����Ua�������	�6�B��Pޗ�����F��%2�L�ղZ��W�q�45�E�]��7#���"��~i�����lAC*QP��/ʵ�h�����~��,�����nU�S���m�j�+�T;�6<�7'��vjE�q®�y:��4,�3��N*�L��ۻ���+o�M�IƉ�M"�y"-n��u�7���b8mv@�����74֚֫Z�����9�D�I��QM� �X._�-���;Ɇ?�=�8Ȇ<c�3Y�&E�/���U퀜���e}�\�P�_5�����>�!௎Or{$	Ad�6���M\�>~�4�$-Yv��+D;��d����*�S��XD�4�Qb��]'��C��z|{KlBa�{����WN����!�?����^��<H$�z�c M����_��`R�t	u𮕉:���̕��q�M�ptL&Q�k��q��vb}z�?�{�D��z�Ba���J{˕*[쌛'��[JF�D���[��ܿe�AX�5�칗
-�:�)�C��e���TEg#�`rj�oY@C��l����u>�!�n!�������)���>m�@� ���$]�������"�V\��U���X��&p�0�JV��zhU]������Vd�49+��I�~�8�{��K��-��V��_H�0��R��vS���	�O{}��"�I�h#tPZ�u���(�;C�,�	R`[7ǣ}^�P$5^rF�E43>�il�����>Yݺ��Ew��¯��\��S�.,�L�9��M&z%���A1�6�HN5����/^�3gx�t&�<ޟ�;¢>�9�pɨ(�\�j ;����v�� Y#&K�Q~o����g`��N�'�v68�/��(��c?���U�m��}��;؀��m���s�U� 0�J%��\�a��F�sə-g�'׽������P��#��<�L$V:���܍���/�<��J�	����.��L��$�me�2. �솸�i̒^�x��}G��kc�rN{*j��д�g������8��r��l��gŚ��z�E���Lo�{W�|��?N8P���"��0�-�౅������
?������..&�+��+E���sYM�*���N���`1���E�33L8��������t|]���e*���ޘ���_Մ\�w�t��.�mR¿�`�a4��J�����xO^G_����T�7��ۺ�e[q1~�L� =
ĸ�9!�u3�oɰ ���Rxb��]�b��:�lF��Ĕ������@n/ωj����JyUxM=� z&�LlC��}|�P���&�40�h�9��B��9��̈c�^�$g`���V�4�e����eY�k�n���O�d�����.M����;)�A����s<���Q�?qZG��`�zpF縷�3ߋ^�;�읕:k�%�e�$b��7��>m� K��6N6W��KP���[Ŭ'�[��]2=
X��rѓ�J�!��U� 'p��p�Nl�hC�a(<'��s:��G����+�ȓ�#݅\�o��h!����U����'��~-����j�Tj^�ġ�!~�����tڲ����T�MM�Y���1�E��6�Qt$���0�A�$��3OE��Q��U�x(o1o �}����r�g]VF��M:�|�M������,_��;���ǹ�@�kߞ,�y��~�򳅬pK���Az,ӼGѮ���]q��Ű>7r���28=�i&}��_��0
$_��9q���N�#�"��e�����8n������
tĚ�O�{�L��g����m�/�B��d�u-��*�-s#Ox�RZ�A��OR`���I�W�z��u�9=g2�b��q��À��"���u�s�C�H��ĕ�w|��G�_ƺ��~Һ�
����V�V�on6���';t�8eg���+oI�O�6�d����r
0���Kk��b @TO�ME?��4Cܞ���XV�:�qRQ�&q"%n�Fy�!+�v�t�afA5�$Ń[����d�H�]�q�3�B���(A����&�S!�� ��H3��!6���(i+�o�峱�ڂ�@�-�:�5oB��(�>q�����=5��f��݃1�BK�>�7������fg�����I�2zt�_�b��t��� S�$u�Joi���U�)�?r}��o����Q�7��G�0{/Eyz��b��XBT_��S}"��;p*�w����h��b���M,5U�`�@S���^��Y�-�3:l�_�l���{[��?�f#2��{�ȭ�����$X	CV)#�Y��}��YZ���6�6I��>a�ƌ�ឿD�o[ٱ�.��6��L{.����O}ʡ�(�H���]+�/*�='5wZY3y�뛋��^��eG�n����MCH�AqM�>,�,3I�X���"9��tt�}����4`Xк�At#VK��R��H���E�}����N�jfѡ�2I�߸�Q/��I'C��ϡ����5�K��'���Ů��Ԕ-�=5{��	���E.�^�������p���z���Z���&���"
nS��r�a�q���B��>Q�&�S�N1��h��,���$�*�-��׆D#����̍���ׄ��,x�7�2����j�&��������~��ʲ�����1�H�99��ΊP���2��sMy�-�>c͈�8}�kAq<����-l8�WV,-ь:$�8��H���(T\5��F9|���9$�vMP-}��U��3X�VKf��GDJ͞�P��^v�JX�5k��cȏo�2�����Ks����ZHߞ3PTړ%EÄ�@3L�����û���l���ͩ���a��M�\�vB�Q<E��r��ac �%Z��j1y�M��ܤ;�-���H͵O��o�����i���CҮ���6Mb�+�(�T#��ٖ�>K��d�s=��RS�GwK����|�:?��~�ׅ	���^	F���{��3���'���w�R�����D�B���<�I�L��Mӭ��R�c���F����Mj3.ڙuf~�6����� "D;Q	~u�l�W��Qn�/���IY�`��j��c����f��#����Τ|�K^(�����/���D�a�E�z����1�G�L�uQ��&t�T?�.@�ER�{��ïS�	LzG�M4���8LCP�?�!���~��e��`6��Vk�o��Qt��\��b�枠U���
�uhT����	YM�Q��U/`��e#?��񆼭�3��D��x�3�dƟ��� �X˖@��a8�����&7��J�6y���|��w�W�dX	5�L�:D��QYЃʵ=�Z��ioq���F�5W���1�[M�X��y�	�zَ�{)� �W�������{�=�6�m��(_��u�Q8݇���e�����������*�ଡ଼G
���!B��kǟ;��22N_�4�65�x�@5.Uu\�j_���\%������	v	��ϼȔB�!��;{c:�W����1{"�xx�"C���R��λ`a�4�&�b����7 �|]�=3��&h.��b��M�`�UĠ� ���h��]JȎu1BI� �v !<��lɁ���[�P�R��A$%T��Af��px�����0�-B��nD�����U����K�r�Ao�Y�ճ�������a�z��O�^*��G�;��OaF�7����P)E�� ���eFq�Ul	hXI�I�=:�@�b'��n5��J2z�q���<��q�b�H��D�#;L-���٦5����F�.�!/����!y�lr[���,��=��}4F_�l�OI�sX��.�n�uRH�gjZ�`F�t���"�i� �6�ס��E�uR�]kQ��\���r��8:KU9�-:�~aw��f��;�C K¢�V�ށG𜌣kH:RbFp�[������)w�d/�[�"�/�l�x ��O`?!�@T�i_Mf3@��&��78ݱ�ز=n��)�N���$:��n�Hk��>≠���'��+�e��Y�/5�yS�?��^�k.o3�BD�F�m��X��{h[bٓŵ�`1\����Yz$�e�a&����.@�tj)�^�Ƨ��6-��qe�(�e,�⪡ъ�d!wk�4+v�6��~ E_�;�j��5�"Y�K3�J50����^~rBS��w廜)F�U(�9}`����I��
�t��wm����
&�^��0������r�o?�
�>��� ���������E
P���w���/�!�L'Yp����_ZNųa��@�H���BCKI��Lz��2�_�r5&I�_sدVjlp�!��ZUKd�7���v�8$�G���r_c�^���O���M�/�H#4<�5oڣ�-.Mt��,�_���2��lo�J���'�	�\�:��?��Z�oS|@܇�4��G���8���6kI�f�����X�8ف��Sse�;%6k���D���}�}�7ˢc:/��'#l�9�pHC!�����y����O/���j`;P���8.�R���ļGb�D���;�~�L,���	��Js"�}����p�8�̕O�d k�LJ"x��n��\�6:�����xx��W"�R�e �c�7'���Cc�Iw�_'�"��'݈�u�I�(����5��z@�4:��8��^����d�	\=>�BY���ts���<<����1m��%�w�\�e3�s211N����S� ���sE��/��&�����8�J�R�)?Jw�q�~������N��Ȗ�2��� Mux ����K���ԗlbX���.Z\�z��!��Q���@&~0�<s����Fʎ��V�ދaVF��J���$��N��^q�PX��a��?
6>�/�Q<�e�KQ a�6���z5��n�D��٧&��7�_f��3I	
�)p/ ��IY:N|(��������$�c�js'����$��l������7SvH�V��ۚ�z���(���7���HfW�n�&�a���.X1��"��4ɷ�ّl=�r�c�����0m�SXq�y3���(y.��eᬓ���A<x��p�EJ�m�Nv�Y�Ǔx��g�-egF��~�7��GNJKx��._���Pђ�%��$��!� ��X?y*��	�W��׋F(�'��߯;�y�����`8)0�j�gȯ�g��p��r0��Q˳���e�����7~ 	�ޑ=� J��_r�zthw��]��~�a%"�6u�PzV_A��rwT�`ﾞ�2/&N��%���љ�,���0n�Cw�WY��b�%�E'C��{�U���y��Y'"��d�<�@@��=^֨RhTE�6��.���㒂;��嘕2�D�����[�]��0������u.��]o�����Y���{G�ƀZ%�����! "ě>�;��3K\*�詌R��Lx�\��G��\B���5A`�"�� �'��~!6 n/����QWo�g�}ʷ~�a�k�'"�dl�=_z�6��e��>��j_kX^I��ë4[E1V3&K��|��Uw���V<6r��[V^�٭�@E��d�J� ��<(��>��싖dk�JdB�~�M�F�f��ϴ��_z���B���Pur�S���pffֻ�ro���k�N_�n�WF*�4;�-�\	ʧJ5X��*��K|s�H�-�\b���8	��1kL^���|�+y~ֵ��7=�Q�j��%�(�3cF�m�9�������Ӝ���yN9�N������U5-�<l���W5�r��)��z+��X�
�DUS�},��s��ʐ�� �.�%vMw��2�'�m��lḳ�x� �̶�[�@$b�3��:vr	�o��I��/4S?l�zA���O��L����6�������4�,�SX@�R�gwo�v�g_�/g���׾�}�o�3�Xۓ��E�]�aO×;��5W,^��#`G��H�j�'J������Ф�H�����B9��bCY�.K��Uo����(Ɗ�
��%c��@ӿ�1VQ�N�ګ�3ယ�X���s��L;p~�2h���?��$��/|��n���[�����٭�����m=�Љ���f��BH~�����-{?�-[��c��6�eT�o(����2/�f�D �&t3��\h�8�n�[��V$��\~8����p�\��yR�ڜ2[�L��.�hH��t�HW��Fy�'պF-ЀYV�-� Yv��a1�T˛oi��2/�T%�1�tTlv�GXeb��5�S���i� �'��}�g�DY��Yj#�x�fI�yI�����ʘ/���� ���O(��YU\�!��J��k�-k�*Z6̹�jǧe�b�?��?��$3w�xÅ��2��xR�x�Fw ƣ�)z�	�2���L�ݛ2�w#�����!x�P%7�n�h5�� ��¶�� ��7X���N`�NZyD��W���ו"B�I��Z�����D�t�EU�6�7�>���P@(��hlB�fe��O�@��)����W�-x���Ӓnwy׬	L�3�ǎ���o���(��+Q$��@mF���8�����g�4�y�M&㨗�H��2��U�<XJ�G��oÑ��Ħ�Qo1L%?�٘�(àNKMea�F�����`.b='�kv�й�o.� K�$Ac��Q�����vm@W���D�Ea䁪��̌�5 ��o�+����Z~初[:�����K�=��q�d^���8���-��΢�NtP@�x��/:0��;R0'��� Gܖ�i��|�����4)��B=��v�ԅ�CYwn�m��;����c[nf��������EQK|Z�FW��vdd�?L�(�o��h܆T���P���5k�A�:���S}�#O�'S��Ƀ1���OU�
X8�أlMI�lo�:򭊶U`��'�b�I[�;/�@GR��\��Ȱ���p�3��v�B?���8���\o�G��|��3Uܙ�v=-�Ď�|����t�\��2���� �f�.vHb��������ؗ9g���>���Pd��-�1g�7R��By�:���:��ӝ�Ζ 	���x�xr~|{tx\���NH`���_����?e%X�c��k.M�@���Ʊ%��ϞT��{'!��%��`�����DNNhƧ��d���/��r�7�k�����E.a�k�|$�B�u����:���$[HΙ��C8Ӧ`D�R!4PA�}�'�����z$�0�^�4�f��A�x��zN�V�D/^0g~o�X�Og����	'�����z�M-����t��p��2�Q��}�ҝ �D��p��A��!SHM�m/V�������P[)������y�)M��N3f׻����b%h�$����V��a��t�W�
�
���5���s�v����䤫{���\�}r�6/�$7��`�֞�ؘ+�����4�HF�KK��(Af��)��B�]��D"qm%�05���Һ����>�A�<J���Vݸ�n���Si�!�����+$]�Bz��'����֤_|0L�	a4-��k*���J>T�a���<9~�UTJYLd���<�z��^���Е6��Q��;������K���o+M��Q��L��8���-��'�th.�U�:���M̉i&Z���i���7k���E~���P^��!��~���Y�>��xz�U� ʴ܁1B�[��H��U��&_���!�H��ԛ�b/�_���IvB����rp�{|��{'���:Ũ8����3u~m��|fY<.XK�F���:X�G����#�H;�CLgiPtãti9nT�p�/�Wo��s�#�������+��/br��c.W��3�����qkZ��6�J��}Z����>��W��ݭ�8�R9��F��I� j���r���o�@k,yӘ�"Z�A�׮�j<Z���
s�����x$����� (6��&ƹ�?C	
�A��Y2�n�����R� MOT�a䐩�?�����g[�� ����
����A���&z����5 $[�ت8�	�>�b$_B��{�h0���6�]����oK�e*��Z6��En-��ʲ׺LosQ��"O�S��S�l=���fܻPu*����i:��0��j�'F���R!�(�W;@lb�f��V=h!}j-)'�r?��
��
)��Ѵ������pG3t���m��ۻ`'r����Y�<t�<AЦr��).��2)N����Õ�=n��|�v�}4�U���ȟ���S�7,4�ZT�'S	1�T�D����l;u�4�x�|9���[�f"@�b'�_����E}�)�w�L�E��R����Ƌ�6����,^RfS�\�Z�鏳�����l6k��Ch�����'<6����C��o�B���qu��j|�5ԅ�3��]�=�I�~�3�gyw�#/o�v9��L��!)f�k�$��������Cn�k#�W8�V��1����\&/p�k��N���M��@�9��5��ݲ0/��`>ŹEq/��_(���j��\`O˭q g0�sib�$��Nl��*����;º�?Yho�����H}�?a
�k"����Dxyٖɯ���mx���9�q]"#I��J�N.�����Y7�@R#���~�K�N�0��}|���XM?N�G,��!
�� ;jf�i��@�So:�8�hQ	Q"nZ�{)�H��C*,���	[�c��t@iuLF\��~\��!<r��i@�}�8mO?#P|�u���d3����?:CR����0O�'������xT����9�X8ƥ�����9n^5m��	�O����9�	*��T�/��Up�W��1��Z�"���-߁�����{��t�nb�&t��/����
�\��5i�8eg�ɔ����	��zYl�Ө=���?NH�L��*y nV�8K�HLȷ����F"F`�����\iq�P�, �71S�6�94j�P����:B<�q��= �(��3J��SC�-��e������H�E�j�&cq�50���A���?���,SL�W&��`�C��O��<c����Z���6��b|HU���/�K�n�)�6�*���W���	>�o����8�ݛۤg�5�	L����%f��϶K&I���`�k�vm��u��� �d��5���p��q,�B�6M��6�T	1!�4��U�� ݙ�Q;���l�đj�@�@�v��o��7�E%�JL�T?�ƙy�p���
8�i�$�!B���R�p4��(d�zN�$�N�TI�{&����n�3o�,�#�1=C	���wf�au�"3f���b��mi��3��k���@9Ϩ����a�;Q��Î�KN��ٞ�\|$�c]P�Q>ڲ���y\�Z��L�D٣�r���wG����:[���J�94y�a?���3�\iQ���I�w��9��1Ǹ�adK�w���k(��)��&�-�����Nc����]Xaw�8��_��R��m�X\Ƣ�1��Q�dn�@p��͔$�}+���U� |	`.�H��6�Z/7���a\H��r���Zzׇ�{��g��y,��2��/U�?k���ף�m����9ԍj� Ah�l:�P��n�FŹ���̹2Q2�Ì��!�X2y�ia&���p�?��&�"�JN�W`'����������o���?��@	:"�����h��u^?T�*�������j� ��d�KߗA-)w������q�؎� �TA���6���x�3l�~�����#|ΟIM� � �a���Z3A&B���١ �fyD�F�`,�̄�1��%��V�CLף�T����=V�xSP���E�֖h�w���ѮM�1aM���`/8���H>���~h����2a��K�5{�k�)h;�Q
2��,eM�密�L�~=��ڎ&U�Wm�%7�I���شI�!�g��R��ug��S�����g����"	%xA���F��Q�y|/˔P��u�@�9b�2'J9jgԺ00_�>�˂��^��$�<������"��B�D�����&�T�����bߵ�������w�}���.z���z~k�%���\#�8U6�x���q����7^/��{�f3�%�m}ėR_x�q=��j���dy�����c��"�HH�~���Ñ�3��S\�W�ۊ�{>���)e9��3����?�Ǡ?Z�oF�}�>�˯�Ŭ���ޘ�: �osJ��0w`F zs$=}�\��q���\�6��LRp7���5j'$Ǻ*����I�|2'^������;��L����#)SoYI�$��F�����s��"��L+���ZO�5�5*�N�g�l�����K �}�I�&9� ����t�)�D�1f§���_LB�W�U�^�x��fn�8�|���']�o�Ar�]%^�ǧe������]$л�4�����g���
͚�^7^"_2Z���timF��r����ː�A��K��Oh��tO�%������������u��ww>�XR�>9����[���w���ke���)2�����ӓ~p�C���U	Yűh�=,n��Fe��򆹤����8iy���Q�~���¹����c!0s�?�s���b͌��d��j7c�fV7S6_���*��r�c_܄]17�.;F��+�֚qU^�Q��
�v��G�hl~XH�o��$?.k�I}�c5�
o�Š�������+�`:R*���lհ��i"�b#瑶Ę�q���z� @FM/1�G�6�_Fp�m���*�wD���-ޱ �����L���\���4D�^�W��N��5ɣ������[<�Q��R��
�
NH �E$�[_�9@�6������D<���H��2�X���'���.Zi��e1��P����(�+rY/YwJ5jx�@������P�l��؋S���$S�+�l���bx_�em#��.g�P��7����8�K���t����'��oP�@�u0��� -ٟ"�U��2`\%���ly�y�0}�PV(k=GW21
r, i�A��ߡp�w؞?�#��-���͂����]����
i�v�/�7nv��sͮ��~���[���<.��vp�ď�~��*=�wqc_����ag&������:���\�K�		9K]^�p�{��Q�}���qv�ؕ���P��B��ۄ$7��
�h����gK������om�g��ME���L�w��6�-2Rv�Z��r����.]=ɖ/����A�+IW�O���
�R,dhL2E�y̾=�C�S)��O�Cc�Rm�����J8<�����Q��7pj:��Ҷ�����������2�����ԟ�����|�z˴=_��Oy��d����`D��a���_c�xδUo�4����\�_ENz3�E�B�Ā���o7M$�ɁC�+��UÏ�$��.R�%� V�� �X����ciU���ٳ�ś|d2Y����m�</ �\v��F����y�[��d#.w��:� ��ͭ�`�k�9�z����&����K"y#̝Ǩ�v}H�rZnq0�"�C�ş��	�y�ȿ�vz�I{+H�g�7$� �F���k�9�`��k��jdWUb���
V�޿�0'r� ~(���l˦xCO�uL���|�0�'��tet���VF+^l�����C��'�6k.�������	f���R�2%����x�L�	*�ɇ�A��0M2ky�ܼ��HF�q���H�=VB����ѕ�EL��Ǳ@h��b �����A`@.��WN{�i��X�C�]�ꝫ�L�L
��Nʼ����rr�67N)^g�8l�����{�x�woU%X�V5���T#�c+����<�f�{�U�ֿi�9(T�@��3q70̳�FA�p"yL�J���-�%x�Z<�>�x̥�if.�TeV��Wr߻%$��k�HUI���c[i#���G�T&3���������u��f���˟��=k�����Re��u�[*�N��PW��?�� LM��s�OWۦ/ڽ�Z�f�o�{���EC\�������"	���k�w�H������j1kc�%��Ğ�W�+�O��E��� ���=g�t�����o_NҒ�4�B�*�l�V���wM$0�3��!P�MBE���þ�f:�;�EM�0����0����
�^��G��M��3p/�)�ǐ+f��j�1*�����2捁oA���t�vw�}�&�$�`������r�V�z$��Ѷ^:V�P��b�Z=���(�v�5G����TsVk�2�T>�%p6~���$��*�y$��R��Q��ǁPF���.y����Ǽ$k�#���bP������8�k��m#������xd�<n�l4�m��V#�t�@�|���<��~�����Ф�7��\�tu�4�7�ww�v�_E=�Q�'��km�
�h���^��∦9�(�7�+ٲ;F��#<�d��"W��i$��^?�&°w��ө\�v�Y4�y�>`������|6�g��]09�>�3��<5a�����H��iO+Ve��tٗ5�7���
�2sG
��#�j �B2 �^#��D��3��5�@�l����/��{��9�Y�ܢ���+��*V��z_jQD?�����Gu���,��I�B�X��X�55��#��a�[]�/j@E9���pfE�󋮕���DZ�+I�j��C�kL��E��SD.�ʖ49���6��i���Z�&���ֹ#q}���×�5�J�N�;Ar��������]ݲ�.�b��H:���c}������(���?�
C3^v:�n�e Z&y���Xl�dd31+̝U�TBʾ@�*�HoG˷v����GE��jRA�h�-��u�;G�������)�$f&��?yŗ	`e?tPk�JK#�J�>�W�W�@���&��8�L}���� A�%x�r�D��)��q�?�g������SsY��Sl����Y�\01v:5^�;�-�5pHa�
^��^u�W����mGEҐ�C�:�� �L��x�@Rյ�ૹȶ�;�7����թ�E�cӐߪ�/��0��:]n�-{O�gD��oY���vs�V�^g�+b�<�8U�T��_b��z�!��6�&j�5�-�p9�b�_�6����"u�(���h�|JQ��-��^����,��WbL�|-V:a֤0�,s��N�"��T��{Ed����X�e� �����sReԄ.���)�_��H^ݖ��M�L^m��^�B-����<�l	�����iSS~n��I>��<�K\�[�;a4��'6�͔*��ҘS��x���"�
 ��ê��Ň�bג=��n]�R�)H.��tK����$'
N���Ξ�7��a�a��y"��-b�>�O2�x<���@�¬�UC�MH+�W�jo1�uK��e"�k �$�`��(l��R�ߥ<����4��F��!0�E<+���2`�uWF_�.(���e7R�'{��p�>�����w8A��sO,����]�������|D7a,[�����-��9�D<���9�B*V�j�rj�mJ@b�D��2N�z�?����<��$�
. ��w(��k�%KiD���f��*�(�i��9�h��s����p��7l6���$&�k�� �l��'�>`����t�->I/3�X�l���X�飻)���~h|��f�DOrV
���	--��,ED3�o���I��sĻ����ZhMY��]�3qs�������i�!�m_��TQ=c�hsC;�Q��=�֩��`�.�M��e�o��vgZ�E���JE>Ȼ	q�Ƅ,�]�fŴ��W��ޑ/MS��V�[+Fc�jG�I8�~��8��i�;,)KWx���6^�v��l鄴�o�u�_�<u���o�c�)euBQ\�U)�ih��~M<�Y։[�7�)��<Y�@D=���w�Ó���n&��(��
�d��b�d�S���z��}�Oo] U�c_B��D��a�"�>2�F��Q-hSЁ	H��sέY�b��-������b���̀��d�6��|q]v�F&/n�eaȖ�CTm�g�ߛ#Z'v��(1~�,��r]Ҍ���<�ǰ=�;AbC���M�oB͜o>��K�a�D�U��e�� h��U�g�Y}�ʞ^�t�H٥l{��YQ_!���:��H�yp�1��J���O=�����fI�w�1U.��1!oZ�S�;�ni)��b?܊�V�A%{�X��s`Kݮ�j[�Lm��Z�� ��i3x����{7�����Rgˤ�d�]��[��K-��J����m�4�r؃2�L�}�M!d���DD:mU7U}��pe��P_�(�4@�O	eJ����R[�_��~��Z�q% ��9��8l	��}e��`�7)��ͥ��|���l=$	�c�=���ȓK���)�o�:���\K��#ğ�[��$h@�z5N��e�A~�kItA�]�f����m�(o��o��~~���1��n-y�W���,�j��d����d����A��|}H�����Y�r��ʢ��>,<?���j0ɣ�6A�p0�^H�7*|���)<�Ř6A�V�GO�J0f��_���zJǅS���Kԭ�a���_(���=�)��`h/���"�&���B�$GʎB����u��Wa��;"wC:�[P��A�b,%���?	����N9W::�ΈjG����,\�ͫ�j��u��
� ��n�ҿB��dieWb�Sq���bu��p�Kj~���QQBӥ%�О_�q!�gr�4�.�6\��苨,�c�yǲ�h7��c�+�7b��?��W~7E��o��9�xaw���/�C�9�@��j�P����D�������?bf��R8�1��_3�.�V�8Z�j %�#�ԍŕ'�e��%��,#�)�g,`����g�y���;�o$��~!��b���f/�h���;â�������P2x���tVJ��	 �dr}����~�y���uK��EY�0x����sL��zr5��Ƞ�p'/7B��͎��]���.�E�R�c�SRh��S���Y�-4�7���|6�ҢL�#�H �,��'ƯLr�u�؄w4�H#�?��瀱ؖrL�)4��vd����F*B䋭�n7~KrmW�jS�"�=�"փ'�������=XJ���4��"o}�G�˛��2��Rr�t&kļ���Ϳ���tg/ߦz�bp$���0E�yI~��؊�S)%�}X1�T���S	QZ����H�KM?O}�W��t�����]�[G�ب@ʁeTײ�I���r�����|�U^�.r�Zbߒ�Ͻ:��͜�CY#�_B�:0��\�m o�f�]���s�гFOpej\J�KM��Ο<K���9��J�ͣ;:2S��8M�r�RZO'�m�۪@�K�j����;��n}jƝZw�&���df"g5��=����,|��̩�fؼa"�˂��q�W��Kh�����T�?�Q���6CZƦ�^{��`�9/�3�*��̀�U��7��ᖲ�|���U�����k)s�Ť��9��[>�u�߲�>���᧾\ŏ�_%�G��Ȇ���o�1�[�AgL!�pI����a� � hR(P�5�>Tɰ~�:��a�w�v+���$�PJ,�V�c��dJÒ\wBΏ�Ѡ�5nn����@�t�J_i�U�GDg��L���X�C�B�I���~Y����}��d�~	Yx�ߔ��[+t�[�nx`�s+�Y>0��׍��7���% *��>$O�v˸�T�;=[}a�����G�L��zD,(�uZYoH;C �<�K�n��.���-�"bBJ��ofH�
�xOM ��;웚��PO�p�F��d`�-���GQ���(
#uے &�i�� <��$�g����x����A.V�ˋwM�g�SE��"�s+�����X,N�z<1C����57�x'�Z�B���<�1� �H?��/>�M�ܻC�%,�#|����|�	�.��|�q�ֈU� =����k������מ��ҬS�2����KY�MI:���T���0�FE��������	B��u�0�U.$����=U�c�ɵ;礨w� �D>�C�G���ʴή�i��zka���[�\��:Ș��>�![�6<�#uz]I�`H�1R�t������3�'+d�ў������5��OEҙu<[VCPS��ܖ�d��'��������G�c��l��I�ٶ�2lY{��~���	'�Hnj�5d	��p^��R���呸A~�:��2�-�ߪ����I`R�URݑ�`~B�֜)���NnԈ��24����;�m[s�͝����N�[���3p��?���IL#�oj*�w��n����14���sE�.53�vI�!���5����n���ɩm��:��?t)a�!5��!(x������3�	M*0}Y���pKZ��Ϻ��0���m��hgD�rߺKq�P"2��^��U��~!��%r�Wh�/��"���h� >s}d,����&oz�?�u���/e��`>�(�;n���y�(5�E��@�LY�M������VO���k��Q�2>�+�v��궈�PBH2�~��B��aO����aͤ�r�h�.]��m�Б��p?���u��a�WT��tSr�u���n��3�s���O(�G�����ߌ����ݖ��V���w���2�xg�SQx��c��u۱�.����J�eFy�6�0��A$>,�L����P4��-#���0�=�lQ��"��_�9k���x[#ӵIM.?�,����;1Qxu���)r�� �tF��l�ɺA'5R�]�udW=�ߤ�@%�?nр��v%=I�B�j�V��!��}`���x���C�P5�=�~��*�"Y<|k/6M��I3���������̩~�M�gm3z�Le1�s��IM�V���U�-yk���f-�����gL2��0釣,/c�J�oGx<����lh WA�	q'p՗;��V�L���iT>29ͨ����3z�K���$��]iv[)��҅'`|��$7�s��л��q{^��6���
濬T�8�Z����&�.U0�4���΁��	����tē�E�!/����je]�����j(���Ze���7�ʾ�c��r~(�.�5얥�I�Uf���6"yf:	Jψ�	���v-�C��L��N,�U-U4'fMQ�Mz�����q�zbM��)T-�\� ��Z��w�4��.mF��^��F���\	�V��!���E�=�'~a���8{���ژS�_�f��}ҵ�EBXM�q�m�� np��,T-#�zyv�A�-��m�^=�M7��f���F��:ꮺ�[�W|~޶e�Ȇ��G7T��{�s90�W���mǠ�"���f����,�d06��`|'��q�Ex���)D��Y-��T ,K�-^,���qN��ʊ�5e�v"��
<�2wL��4����Ի��ES��(�N�������+�*.��U'�1�J�|ɥ��d��^���2�! �\�O׀	~��o;>������/��%M���{�A
���:U��/�%]D��i������j΄��%7�l�gt@�nK�-�������m��i���kw{$d1�5�S^;彞�$4��꾐����<������w�|�r±v>��I��^M���xr�A�zE�dm����w��&G��b0)e��J�5J��K��^*��ɤ@b�176[8J���-�/y�����'���I*��U=%�E�cA�7`�+ó������X���{Ց�G�פؾ��>��2�B`���A*fg%\�C�(�ԣU��N}����@��A+��`_U.�V��(f5ncʟ+.��~�a�y��<�D�ZK��򵮖֙�u�6�ΒZ>z��X�7�W�n��(�&�$���^B>Yd�cxC�{�$ON��"y�/]z3�J����6��w��6��`�T+��=�S�X�s+��A�����-q*����y�fۑ��K}�l��2������~Ʒ��l5{�oό���<fc"��w����J|nʜT���L��|��iR$9�><2��c�*�2��xg���_���t"X�U4��+�k�ImN�Q�Fş/5��_��H2��k�}���s�z'��<����^q<h��A�df���0 �r���<��n��Mck�9�a{l�F��.���#b�lZ�f��y:���0Kl�9
�M�뤉O\H@�R��f�C�V�r����(���dhU��SA���5��6��Y[��?u��D9o��h����<�bԩ>���5q�x�M��b�Mw�lY�K&l�k!c�B�@�f�K꠩U�j��}S��'��\֘-�y<To��U�Q������ϻ�:����
��j^���[R��D-aSw��q^��o�V�p�J��	;���I7;��ls�ŵ��GW׽�2����� ��<w���Y�v!�ޏ���f������I5�و�>t�6�PY^�ˬ���xU 7��H�fA��,2���s���@�]�EER�'�*T*mh�G�SvKH��@���jzS{����r�J0҃o1�Q��NJIiS�H&���v�#i����4���K�*��I0�����cűֶ��r"�{	�:�q���x�� ���š9</(5��Mx��=fyX"��j�A6��ve�%."j��d+��44��#�[l��z���-��22�񖧙/�1��'eX4�/�6|��1�<����ˮ�&"u,�f������p�c�/)��TA;��~v���V�m5�ua��\%��0V��7T��T>�Ua�K���B���8��d�V�t�[j�Vg b�rSu�%=MCG��CҪ����	:9��O
�%L�`�~p����v�̊��y���\=��f�hO1�:I�q��gBW�<�t�=�4V�t��.���)�V�-�:�U�2�FYGm�~JT��i���.|�������#=��Y� P��`M<E\�\�x��x�����+���'aI�Z�ura��f��}ĹZd*�#�t1=�+��4x�a�v�9#&��a�b��;aVcfڙ�p���8�3P�>M��^�)tX�c���S��'$���괦��?�;R�]3�P񴸸��MBX�5�PPs4��HC|q�L���U��Hg�ڑ�E�3T��8�?�s>2l"Q$���z�b��u M�Mh�$�T�c��4���N�b���Uoo��vv I�l�����9?��>���!KBY���c<
�U�<y>���>�G��Z��2z�E\t��G�{��F�=�u��+�D��o�۽�.�\���+la5w����FٳE;�NY�~+�Q��<��k�{�j2|R?�md�3�����h�k|"\+(�/��4�N�,{W�#;oc���ĳ�t=��`5,e�al{qìXF���McY ���$4g~��
�H9h8���.��(VG��|�.8wAa�}�W��y��!�k'��&d�:�VB���@H��#����l8�$�4����	�
jy6�_��k>����( h�)]l�!|9�n�\v}�� �/���{Z��u~��������gd,QbD���q�*1r�A��A4��:�ү���Ԯ�!{�]v#x>���,��G־)(KW�(ĆJ۴Ւ_ ;Q�0@,�� ���h�L��E�$�܊�쬝�wI�_T�wi"���$�)�[8�N?}+{̝t,����̒���j+�(g����,+'�-��X�?����ɯ�2�؞}��΋������T�I0�I�Z5ɍ;n�Tx?'S3BQb�Q��� ��l5H��\R��w6�а�ެ�|W��sO7���A��&D3��Aa_ ;��HĞM�e�dWѾ��}�S��"���1(K}=�8�K>r����jM4d�����3�H���PX���aM5~�X������� ��?���Twug��fe	&S(ɒf�9����A�f�Jќu�Q��<!��=l��I�B��T��fZ(z�H�f�c��y5'6������L�Sx��>(I+���+Hǳ�u�?z��1�p0��C�}Ͳ_¬���喍O-���Y��'�|4�Y�����:�p�:#'��Js��Q�[MXWA����xo�R�y*y��({#%h(������zg�ͨ4jV��c�����1� �h�t����SZ6T_�i K֬��`����		�`�\�^2T�J(9"�o�RϚ��M�����V �D�E������gW"d�@�T�ˇH�c��e�O���M	��C�`�D��Y���6���{Jѫ�]D)x2���uEk:Щ��#zԳ��kK��b_��Ra���{kv���o�8o�fE1�h5�\��-D1�	�/�����3��T�\�~�"�_�s�^�lr��i�
>�MS'��(��!v$�H^�Qk�ʞ0:�)�ڬ���5X/�at�୳v�z^S��:��t�B{_��^q1�mdLPi=pV�g������!qx�g�p+2�^.W����~�A����%�N�F����r~cX�Եu��{ߘ��� )�i�ӝl�9�P�m��������{DL�˽B�}����9�T����^�QMaD�ʶ�
�s��86�[�U�RƠΈX�3E"��Մ�s��o��A3թ
�XѼ�K��Jf4�C�x�����^�5��  �_-�[�ɩ��i��)w�;��pOxA�BVI��{/����0�?���|��_�q�`g+��Y���q��Y�Fx�}�0B�i�Fj����1t��zT�ޯ2�0��cH�j�q���T�Ox�#�l�?�8x��BC5�]�����l�N��T��\59�MV�.|RL M�d��6�
���3.��j���b���i�/b�0 �61� ���$q��ߪ�}%��pR��"!��M�
NBm
Jl�k�կ�M=�[�LK�ڎ�)��/D�����C"mW!���6E����B��n���3�S`Po`�¥�G�\ ������A �~٩j��J佨!rKí�Q�|��v�o�+����l������F��T�;J�'>�����o��v�����e�,I��ϸZ05��A��E�%
٘���P�4����o�oV��2�l:�&N�D���JA�a�� r�|��(��o��eM./񡜐�����,G}4��_�2���֎ v�à{l���@��P;���R��2����!�hH��L���$Z����q�V�^ i�y�C	Д���b��3�/\U�z�l���R��Lb�3o�cᦺ�r���+���p1UW+���/�ԑݏ�:F�79��:�?-��
#Av-�+����"��-T��(���	,u��ȴ��Ľ�ÿ�:�1�v�f?P���S��p�î+y�	/P��_g�~�.�]��_>��KKs�O �`6��Ld����&��	�DˑV�$����'E=6'����g'XJ����;�R�#Mv�đ�(���(AvbX5f�=O�+0�E~����i�`�R���'�N��:yB�L�'���fB�M���H��m(6��iL�9Y�H��-B��t��;OS{B�G�cT<g
G��C<o�mX����//���G&��b�p�Os�oɀ�}��W�B�	x*�4��H"�u�r	1����x����'�1P�s��Ǡ�}�Q�����,f���寎���aC�=9����8��D��l۽	ɟ��)##���=j)�=�߹��A��*�-B2�,}J8��pPdZ��������7�����^t�C%�/o�M�(�"MF[n��ݶ_��4�����|ݻ�r#��*�L��]�8(p/=�C�&��(;�j�db<�9z�����臬��8,߰�n/L�������Hu��J�o�CY���J����-��S'�l��#�浸a+>�9ȗ��L�?7�s�i��R�$pd��B���^I�yX5�'��(�e���y���N۷[s�,0�P��{{���Am�a����0l�
;����=�DC<�V[w-3�aO��p;�����&	�S��吹a���+Q�����=��ɚ�fꂡ��zzੲ[�о����9b0�s��T�:����nJ\"�֍(T9�l�_\ƭ�V�Pl�F\�B�\�)�&�:��WNF����JR���t�L�ݧkR�GK���H/I,������TS+���`�*"�çK������l7y�h�@�OE��W5b��"���9��N��3���ͫk�.ab���K/OG�X�^v��x�Qە�&'�N��(��?.R''�y��&y6�����(�}��x=Op�/d&��	�x71\Cw����>�Ee&��"��#%�Ƹ���"q �y�vU��ߋ���4�	_ҔbRy�M�n���ϩ'��/��L-?��S3�]�nr r�6l��be���S�L�U*�t�Z�{Ke/9��Y�(W�&W"��v4QZ�P����B�%������KhVv�_�0�<&�������`�r?�T��7a�����P��j����7�A���-ކi����ß:�
���CI��l���誰ܩKV6m55p�
��{A�I���H*�A���C������gtB�I����-؍$IfEJO��T�*�B�T���Jb��� 3H�[��d�ּ^`��Pp�E���b��ͺ�����n�,C��}*=m͑T�c��H�ۢ����3�pQ2��$���vF����:����:7Z����j�hH��ߥ�c0���ȀÚ��:JK�W@n(�_��)މ����� 6��g����W�TC�!e_i��ԑ�vZٓwo{T�yp�C���L��Ez�������ZB5�����Y�+{:��:���<*�vV�q���,6�7V��\[K��KW��P��t��1�F��<�S��hq*�Խ��7��N:���|�l�ʖ���|MA1eXB�y;�����18��w�z��z}1^�GZ>�ZU��π���m4��G�8���ᥟ����_v�'����qF��/���2�k��@P�;�SW뾛��c�S�:��ּ��Fi�F�X�W|`�M��c(��8�&�=���T�	�y�A˷+�;����P8�ƕcr�P����mfK��g�r�sF����zT�'>��:5ȧͮ�_���Ð���;��w�W��Է4@�;��nY�\V�Bm���s�$�sQ4����A��8[�V���[Kz��͂��m�	@WN��}|S\�ׂn&�H;Wg����i`�Z�c�]��宝�7��Ά�R��t�ڒ�7�eX�ide��V+�$P�ټČ�;�b��\�}]�m�ծ�qи��tSzuNa$�[���Jg&�4�D��/+�wM��G�ŦX�]`��9��ց���7�wi����9����q�~!j��/-�\�Z�>�� �6c�`�e�g�TA��I�{�ev���c�2�J�r����z�ǭuYߛ��J��&�q.LcRU���.[�6���]�0��{���+�1Z��®�B�_f�/�
y	9�uy�T�S�%w�!��V^�\P+fAA����I�j����C^�u��l��׷Ǉy���%ٿ.�x�@���	�ׇM��#��Jv5��׌��oH��K`�z���W�X��H����w0�6�{�3�2���$�u{Iس��!�e�^�7n�H���2R��NW��B����L0|�rt�sj�|&#�{M�S_�ǂ[�Zp�I19�/�C�7IXq��)s�'���<@Y�ƍ�������Kc BM����G��� ��hb��P`���Yp��A���.������V���^�2�;o@[,� ϫ����jx�O,u����4�?�B�H�3@×��_�p���v@s_恐"�ӻvuy6�d�7�&�<u5pIPa=���3y^=eDK����C��#�o��:�P��Y��O����.�53� �!����뱪���`	� ̅�z�y��I�cP#K+�F��<}o����H�x����.8��lq�}���1�9!��W��x/�M��3x�`�����_�����ѩ^iJJP���ɤ��-yk�4X��>�L�
ӗV�>�KH�(ص�W�1���@��G� ?���������ܴ�9���E�o26�� !6�si�t��]y*b�:Ԭ��OfY*�cu���y�cMm���j�?�ĝ�e.�mز{��l���Ҡ#^TZߺ6r�����+����)kПv�+T��r���e�*��*�1<�q|-z�`�#�[�����c̊���m���F�0fҗ�>�D���Om>hmq�����p�J+F?���dPnΚ��;"������)_p��"���0a�{���%���2*A��	i�f�^���I�������:y�l�P��'��oai��-�k����I_�����r��(5��������n�)�u	X$��՝KUh�y��n��p2d�����e�M{��^�3������jP�c��w��.[��0#_��y꒮���U��܇��� �����
�߇䵼�Э�>G'�;��`k�X�=�4c5t�/j��Y�����r�����<{%N��1M� ND��H�y�U?tCv7����p��C!��|ce�;U��������}_�$)\��{rX~f:�Z��`���&{�z��^�ʟ3&�Ԩ�,p�h��y��@F�?��Zp��eni�F�.�fF�&�z~�F�dZ�t͵ק�M��jZ/#մ�9����Z�ʃ��߀�Uy5�">X7e��r���O�(,� �)Q�G�A�����FsB��A�w��Ѵ� dJ?���3���p�Ԙ������"ΊF4p�B��� ������Y5�2lÄ�}��|	�!�	��
�m�����B�=:����k�8x��E�c�N�;�7+�J�x�ԟ]B@�R���F1FfYS�r��BlK�)_�O�Ɛ�x���0�U�p	7�V	��::��X.ϓ��w�=U��
��-X ;�(���?��ba��A��s��Ɵ-o��[���c��DVkik~K�b�W����Xoˋs3�b{E���t�:�%eV_��|�����Z�vZ5E�_Bࢡ}[�I���N�kM�(��}B�`�s�Hc��T��+~�BVwy�$��5c��C�JŔ7�$��Oe^_�-�+Ґx.��^ �;Խ�
9�I�t���ʵg"��@�OVn�ֽzׇ��D�<C,+��66��r\7�TDTp\�����R����e�܁�u��XsU�+�R�9�'"��ב��f�Ī�:�T���8[�;�#�˫� j��j�ʔ�I<�ynG\z��00�,uۮ�]e�C��^�(Ԍ`U&�9 �vM'�Vm�����^!s����_�����Ez���#��d9�rt�e�4��- i����<A�� =ļ�NG�I��/�p��u%�ԅR����WjZ��� ��k�i��?2�8qDM�������Ҳ�']������2�9.zOt���V�׽�~�l>u�����di�y���n�L3mj�U��c�'����I�p����L������#N[�F��n���qfMz�cb2f��F`��t����C\։�هd\��E�ʱ�B��E֜' ���/�3Z����ކ#����C�Y�Uau�B?��׶W� &�R����(_��d�F�K��+�7vq#�b���/Z��Q��]L�̔�F�	a������?Lqk!v���.�<R�\о���g�WW�B�%�a�<�1��������HA�U	��F�N�eAN������뚚�W�^t����&hw���x��n��[��D���EH��T��E A�u�$�Z�+J,C��pyT�
�?Y��������=O�8�Fb� x�(�8�b�q�b���$�}����{W�ԶG��������@l�og���s{��G~'h��z������$��d�j�e��[l��;}�����#π�{|2۹_�g(Կn|iQ���Q1�e��������౭��$Ƙn��"b�ys��*>z��#�V1�/�+�wy��5$�_84�|Y�f��M;F�|q���T2^Q�u�5� A�V_�_?F�j*�ÃY�s����W� m�e��RL�3�Q����-δ��2�����>�%xg��fCYra��Z������ ��Y �XE��������t����h��F�v�Ш���4bu��b������g1�����M� Ŏ��P�YD�"\��|�������[4ygQÀ~�]��R�߸�U�z���Q|��1_�,�t9��7e�7�H�������~���³�O�@8�6V^���M����d�����ga�� Oj��(
xɨF����g���|�~��<(y�m��:��lZR�]4�QB��֠��*�(�7���ea=�@�����ޕ���L���Je��adE=��ǥV(8V��#�T$"��x̿�W5f�s!ȅ��Φ�-�j��6O��w�(�s��R�($�s٭� yl�Z���i&�mO9���DI�Q#X������'�1���1�#J}��<�3�um��:�V���L������vOv�(��.�b�/y��4�H ��Q|�P�|7֝�sY�j6T�m�3'�fj.�������<Q�i%\dr$��ֲLI�r �,�(Xt�`�3�L��k9�%j�j�NB��&��`G�_/�WG�ZR<f[���]7󍍭�mw�G�<��#،
M�z0k�͑Ż��7��'�-�`/��+&O� n� U�"������yL��TE�-�S~���YZtS�Vy���0c\��
�ꍔ܏ky�s��:c'F��VBzV�^�w~c��)��k>�	�~*�E�01��0�>'��a�HCg�=b��QJ�	�j�Pp�oZQ�nJ������u��X��Ԃ%��7��-g78�,7h�r�X�>&l0�ή�
�3l�����?�=��^�jv��KP��Mw�I��l.�0�Q���l���G9�s
�6y���8�&�l��
�1�um)��q(���Ǚ �гNE�خ�X�\5k�}(4�(]�ֶi@��S|#��&��\{pl@�����0�zp�G��$cF'BR,Ć�wO������D]��W�S��FJ��
z��3[=�n�/7��n���P/s��"WI�/y-'3x�<�ys̷�6�vD��"B�w3�M]8�9�����Z��apX������x��վ�%�&l��\�4���y�J������5t��!�.���f��=� =GF� iU��vE%�E�lB�M�t��q��t��B蔱{�g]�1�
ͼ�<��d/�1i3o:-~�Ko:ev��:wS�hV�r������1�m���/�c��&���D���95��ElS'�S���㥞��~d�yUN+h�3r�0l�	&��N�
��D�Qy!#Zs�c�p�К`�/i�f�`l]Wm�,aH�?7��4!	�y�Z�? h��cЍ[�:ه���I^�,���z���>�;�n��fd=U!xs^5���4o)5cݕ�ܱ�j�������?�"-��T�b�IX>?<y)�
�{vz�p=΃���5TrC�Sb&�>�-��_��ޭD�DO���
<�J���Y�8K���/�z~��}@�n�1�J�܉ �ӹ�Z��(��=HR0�'D��&=O�~�BM搐��x���i4���?�6{%�_���+�R�����P�W	=4T�u�Qg�q��EC{�!|��ԯNmGL�r|�*�Q��M���΄�<�g�~�7!O��BU4"�->�>�}��J{O�(#w#P��ԦV��r��Q&�]\-͘	�7�Px-��0��q���4��:�=~�bN`"�De�� ���z��),�^��EZ��Q�z��uG҉�[q/���wڈ&�=^ �ǧ�Y��P��c,�OR���b�f��mGW�*�E ?	�t"�:x�|%ߺ��E`�q��]�F���z��� ��{� Х�e�T�lMHM�T	)���zE����@�8��@�)� m��K� ����'�@m��CT���绀��.�r��x!�/�.�{��)�.�=��M�
ؖ�T�/��;���{ն���wy�v�݂��$L��)�K3��|$���P�<>Q��H
���!-_���>L�sؚ��L�8�?,�|�~�{�;��6��5y���+P�R5���t�2���e}H��5��� ��K���YZ�9Y�bB�q�<��ɇO7ϑ�m��5�!A&��G"1"[$��i�p�R�� >����9bv#'�J���֓s�6ʟ���V�a�2mp*����'faG�bl`b�O)���)��b��@4�/x�E,F���!�U���|$Mϱ0�'�;o�f���?�d4��"Wڬ�/Oz�v3Ӯo�
W�F���u��lwHwo]�=�]���=>���XF;��U�%&��{-���]v|��4¾\|���3�Ǳ��7F���g��Z}d�-ԼI<ܮ�	=d�re������t�����T�do^+)�k�6��:n����J����`O���9�b6h��)�� ��O��~�����v��5 ��ۍ��R;��X�3�~�����6�<Vmg&y�3�/XK߼[�����Z/�(%��X֐�XQ	w���TE2#�����k���{�'�ա��𢒾F��  |���ÀY���A�:��f�z�v5�!�[�4�p�6�Y(�5�����< Ơ�B�7%J���;��S���g�RXu�t���7�n��0�Q6�O�8�k/�ܡɂB2�B-��0NE-�p�)$�\�y7n�rn`kU@Ճ��5d}�K�������bn�����j�MC����7��.����*�' uEl�}\�I.C��p@��n��=ײ9��x�[Q.��~5�Pɜܗ�:ԣ�7��=?FN�%oK<ɖh�sp�p����p��ȝY�V���:o��HE��ӷ�|����~�Ω:�D�ZM��96�Ə)S��ϸR�>�:�7P\�aӶ稤"�����&�6cRB��� �Sc쐲��]ϵ]̗��5Q,�Բd�2jM��7Pb�y�-��j�+K��;�]t��>�%p%�Y�]N2�eы9Sy����Kx�TD3�����I7�#�S�ywhQg��������$=�- ���nq�^{]��d�g ���s�]������0�f��U��mz���u������K��}�}��l����
$����*�Vn
���.'������M����F�2f�8����-��˱ly�B�D͚i�]U�D���$��[9��>ʶg�q�3(���A�a*�!�	��6���7!�2��5!�/>`>;��ǜ "��<zec~���ú� :w�dϩ��Y�e�73v��>:��\<���fj6���z�L��q֐�QHs��ɇ/���6*���,g���kk���}Pv=���aHJ	��2�e=fh�1"���?�)���H݋x��@�������ܠx8QѽQ�;�Bߟ)�G��8^��IE�re�c�u�2]�=�"St�V�;8@ � �����,>:p��Y�	���8"�WF�I�㰐�;a�y 	XE�/��]���z����^����H�2��b�d���x�=��Ar\��T*ψ��қ���\ h$���0<�������(�0����<O�'8H=�p��N��4��?�^jB��C�0�<���z�����к���P�H8f1�=�5'af�M���~���|d��b���Z��P��,���;?���+�d�D�F<}�C�C��7�D��FW�a�&J�3�ٚ��{c�B_��~f��艟6�$4�����<9����(��
�ofT!�hq�,W&޳�ڨ�+����\�<;�(�Ǆ�-T1f9qzT�/4�)����#�9_��/���r�� �?e���Ѭ��jz�$�]>��}:�dO�p���"P5�z(f����.��;���úEB��<��Fj�$�����tK�k�6�)̰�1�|������͕��7UN��H���CL'��Dp�BVP��Y�^h��3��x�b]���p�g��T����V{2�JF^�Ef���v\G�?�m�W �Yn�x��6z�[>RCc0B�J�!Y���(,{�<N�e��;�[{�Ǥ���}�XC�2F�㶮�(��Z �攘5���l�@3Q���x4۶il��s{J�lU V���6OOWR'���-��h�y`��qc��*��ݑ��=ZW'��ǉ��n�s��c��1��T���Z�$a8��.K��Z�p�rB,DXԎN`i������27��$��h�M��ػ���}����d�����V2dX����9�(Ź!�N�g�O�m��T��C�c&�0j_�QK��یGSm��#	��h`�T�4	,3"k2�c�)����s���@��P�4[��
|#�P��|���uF��|8�<���l���e�R�G1��*���	��pђ��x��-�4v՜�2̝�y	��n��+�3���A{���?�Q�?/:NtP������"fT&��v?ߡ-�k�>G�Q��W+JS;W��Hk�C�l��Z�����GI�6�rlªYPʠ��'�肘7��T��3/K����ۯң�c�v�Ne<�̑�Z���6���yihp��~����G1k%@k�$�0��Tr�?�K#�K7���;)�u�&�Qh���Sz��C2;�T��̊iͽI��я.��{u��hR��T�f��N~d.�Q��A9�v>���̬�t�'��쨵[i���j��"­�m��~,�;c~K捽�2x7��vfG�)\���H-%&�n�j������T�D�����%�lM]'aٷ�S]�c셑˝ͧ��:�TX��y� -�C3O�	~��O���%*8�<Q�O����q�̙��?�ޅ���U�&э�|�mݶ������74wh�p�56�>8���k��4�Uj�4��JK�y{�ō�xFGFSks3��/�V���Ѓ a���"�
�L��#����a��iT�V荾�m��-0���c,���ۀ���[�����*u�nt�έ���~�?��h��^�~���OS�zwp�A4zl�!MJս\�%(Ϡ^�_ƈ^f���,s"�v3;�-e�-���Iy�Nni*'2��d�͡��c�gT�#�Y��~;|� )��x��Բ�3�85�ϴ�i
����������!��$�h�~QrY&����W0�v�Ơ�ԮeC���������E�(���GP-g��`Jq��<���5oQ��v�e?4�f����l���zB��%ŵ���39//6�Q0VB�_JA�Å���J�t�f����>��+Ǩcޣ�Z�[�O��i�a���E=q�	��`����9��p���E�l�`��:�ػ{��S;-��o5n|�zYx�{�z�i�:��i0��.ɏ��J����g�K���##w�b����	|���!tH̐��s���������$6��3)_i���S<C7���#���ܯ��l�I.�'���V�3F
����H2��⊶�w��!,�l�N��a:.�{�÷�_-��F��7}��-1�>����ь�B<�`��&�xw�&�΀@5�&O_b��}�rn3}f$S�!�!�áq4�k�<UJ�������� �4��F���.��ڋ��_���o� "s�������<� ;Q��W.�0vI&����m�iN>�#3l��-]���5�
��:(�����J{��#�b�yX�cU�A�ʌ����.�J�z�?�q��;����!�@�Pp�s��3�g� M���Kɹ���"O��xA�a���^�I�]�p�j��Ԩ�K���QA9�����0��,���\^M��,N�`���y\��S�9��/��N�[D��IS��;ߗ?�Lh(,��;��_����b݉�;$fM�A=�uA�:�hC&To�=z�D����qMxh������]�
���y�yT�Y<�)l��� }��/�:.JH(����l�	T7��zp���	5kO�sO8�t6�"�ad�EJ����P�A�39���YȖ�ɵ��9М��MN�|SZ}5�f�/�#(gR@�m��ZЀn3rA�c�q��vU�O}��;�ke�#�6iX�������f�r�V*9�����2w�����5�P��%�#g޸)�EӶ<Ɵr��~˸��Y��t+T��Kު��|L���܌Ic)s�Ⱦ2��o��m�'����D��]��yT�<W�7/� Q¸,%�c~�E�J��� �uA��M-󥋫����u�n<@[�u9!�.�@T[��6ED�/Y��;�$��d���Č��$�B���\ڰ���+�<��yV�wa�
)�п��Ca�7�\����.��v�	��k	Fk��t�p=�h�+��I���\�Ƣ�I�& �s'"y0�g���V��b3��v�Zg��A��!^u��`EW��JL��Yf��M�쨮fD4�,�(x?�����;/��Fa�eU�A�s�2��e��a���JSM�ޢzU��$��[+�q��j�2+En79���&S���C�)�T�����sy��wB�����x�陲,E��{\6�l.R+
�D,ò��}��]*����Q�l<��-B�q�f+w��* �
�/���F�C=�%~灅(Ϗ)i~s���|����H��4�l.=����9F��������bl\�Y<���~��
̯�-��o��)�S�"{f�K9	 ��!��z���+��i(�F�j֦F6���@���1ǰݼ�1jЙ�te�"� �d�����97���u��!gkdƺ�{K[_u��%*
��g>���}�0�|7�K��?<��.$xp&����������"	�2zqz�~�l��佂^�0�����%K\�̺�M���ڜ��W��+v'65���b �я�rb~p=�����۴��L�=^��zmh�&��YB�D��m]����u"�oh;=��&F�>�P��|$4�x��Cww���$�ң;���9��/�ؑ�����a���MD��ڳ�j/��g+\�]�&5��͌$�gץ�n�����zR�L?w
������sQ�W�"���5�	f�]�����Q���x�c�����i��r*�Tx$X�W6�$D�@�P�+b
Vy�����m�I�S�@P�h�	`����DH�~L;�=��+�������(v�y {�٥�Dpr���2
'	����C<jf�g�1���T����+q�vR��v I�lQ�&�{+��;}<�t�E�xUVm�	]���'��#����	s�X��<U��{�r����WM���0=��u��MF�ς��IX��ǝȯ��	�ЖWgh��K-Ž�֌N�k?$�Y���}k�^v��%Q��Y`6Y��p��iłG�;|���S�F����w�o₂�{KH�QO(SF��x��G��a�2P�I��x)S��e%��[��<�j�$���4O;�>�h�nF'�}����;3��Ngⷹ��
/�1!��oN�Z ��v�k2,.y�ǽ`T�H���8�R��-B=���rFԛ&"��;'�1�@�G���f��֊BF_�}p���V�?�U����Wk��r@��)�];�L<��$��`�4#����&�K��k5�)��9v!�0��+.�,('݈�����M�d{M���u��N�����Dyz�k�HOz�ֽ��&��
��cD���d��;<!�X�t���])O7�P[��sj!b��b����j��c�	���J��aK�!�k2W{G��Vz	�Փ?�%����Q���\�ɹk��1:k�m�X����x62�$h>�V%�ë�<�y�AX0�u�6U��k���͗h� ��\A�G1�W���VG�s	Ԉ�����������͛������/X��*��5�������iR��#�͞�;I��)e�8[��5���+|���� 	��y�A6����:<���v�-K�M���F~CV-���~8ZJ�$��HZ�y�=)X�o`�Z�Mq+!7�g�B��pF���;�_Ms�{�<&:�:�NF@Wӽ�L$�(�ʄo0��n�+�匌�AЍ�X�5r�5b]et��Sf ��4�
NA,#Ω���p+�J��c@���~���ȳ�̟Y���˙�|��9�G����u�X��%f7��ݷ�P)�g����gr�"W0��_����E-��N�Å�� Q�_���0���u=(��
�����&\�pll(�p�傿-o�/�2�/0q�R�ׄW�`|�	cW�l`�a�C�T�&��8�
��I��Gծb�l�l�gQ��J�`�58"�$�)st�:���Ǯ�,`�E�o)̉�g}��C�l:E�RM�,��%��΄�O�y �HZ�;��t���"�4.J\�Υ� }ݯ6�ڙ{ ��Q�]��� �%dz��qWQ��'�8j�
�Шt�����RO�k��s��?~k3T���H�&)�_��;6%SG ���e��7F
e�9'	�N{�9�3y�6�n'?�6։
p�GG��	��d{���I=%Ce�g�V����f/��_8D���ޝ�|���
����[���q�����I���uf8ɽ��V7y����f6c��ۘ�Ga���'�On��S�8��V+�A��0�Ę�S�[^u���}7A���;&#�q��8���u���Q�_��R��ҵD�3V�7(o�� �k	Sf��Y(��I��6h�s/e�Ju�l(K���lMN���%Ы�����ܑ��A�8�Gi��$c�wc5��Bg���To�d"�y��ⴱ��1��%z�5P5��D�?c��V�(z��74&?Y��v�K�?L�1�b�8[W�S�v�Z�t�B�O��r��aMi$��D��i^r>��d)l�����N��S����9.G�D�v.����S�#���ǉJ������붽��MC�BH"�itP	DdwS�}c��Vۭ�RE��<�^Kx�p�֯pQ��E�O�W,���Ŧ�]�pFn��>�c�_��A�5�0Po�1�y��~�^q�sN�M��A�ŋ-U�6ǎ��\���H���AzJmO�M���|i��0l��"�U=g�N��,�V�o1��ua��~�[�'Ҵ��&��c}3Oz�hu|� �r�@�Ӽ���v-�m�fDiO%��z��7,}�	*���n��ʜ1E��AE�����sw���������izĩ�����z��W=H����Ul] ��0����m]�>�x�G�!�:kь[�_u����X���~W���A�K��fhǬ�2n<EYE����j���ޚ�TY��:!L�eVt�ϲ��A��Q�:��DG�&G��Ê؅�nq,C���:�Mc���[�J�QlF�1��}�Y�ى[5o�7N��/�Z�V]�-1ۭ�y�D�;<U�;S�E�1�� -�J���o��FQ '�1�Dۯ <�������Ip"uP�9�"�J�~�Q�.��_�Mc���o�ݜ���ض�V���	+��qݎ����֌�#@��$��;��<���@@�t^.�Vk��b�v>AXn��������}}�v�15��Skr�5���iyV�_���^5��H����b4����N��6�dFdoL88��7�I�	�T��gf*ۊ#�v?��U����8m�t��F�^K*�;��{&
�u�`	���u����U�:L?�{v�r���A4�2\��{[�(�Ӊc��7�X�:���'���~.h����%�68���{\ke�`��� �S�p�γ��Q)F�;�y�!Q�����ع%��7��i�i�.C�+ջ���h��A��Z����KF'.�t�t�yx��
)�g^4C����H��0b��٠۝O�M۰r�6G�N��O����n�+rEޕ+�Њ����H�`c��	�zq65���n���F�b�~�0���9���n�]��Fpm��r�o�ö���f�����n]!<:RSE�7��� �,鰵ͲQ�|>Q��F��Ъ~���躁�#o��<���B��g^���fދ���<�*Q�w��c������]
er3"Nzt���;�vJ:_�b�_�����ZqKM/�`XA>7�1CȽ����ň��<�Ki൸�a�Z����!$\�=}L�Ƌ!�9N���g^�3C�&3��{���@���Z�)�9�S����1�B썢r��k>��ݲ�6�}�^)U�Ю����E���yR~izy���pi�Q\\ؕ�� ��G�Z�iH���Y�n�#�:C{2c�-�BD9�ͯ�����oFk��(b5#6�.嬪��a~���&c�l��L�1+���"A�Z��z�S��\�Tb�G���:u�p��6c��і�>� /��P�'�B���eM���S�Qe�5�=�I{�|�)$�b���g|c$/�^iƤ>M�r���5J_�an�!7�{��ᚒ��MZ3��u]ӭ�����>V�c��O��|�*:*W�keB���z)*�>b�8��|/������͟-Q<7�+G3�ɚ��g�+a�+v�AA���!��R��\	�呂��ӓ���_��?��K:���˿`)���m��P沍�`)�-x ٓ�d.q�o�^��3�k0�;)=I{z��a���T���}�͞I�K�Y�I�����p�r� ��z��%�9��ѼZ7����n�|��~�+  �9S��:>��COF#�
B��o�_1#%��AϿd�E��z�?}ÕZ�j_`5X����/�`HJ˻�m�G5����QM��d�Z����_�[��w.�-� h4���fa�#9�o���|.��SM�qr�p�Zw���KfS>(���6�Z���z����oz���8����Wp�hzn��o&�@�3+|��ҧ?%��h��be~�H*���>1�ϚŕJ�R�����r��U�":��e������:��{�N���S�
����g���Q�Q9n��ゝD��gK'�IUw��ytfK%:��)C���L�]��m���v��~��e��E��?C��4��f�f���A8���4�E�	&�o���\��S�I�ٶ�S[|`7���uӎ�j�����JZAh��Zw�{%����M��Jہ1�=K���aTb�]�@�
Gp��_�6?��Df�6 �'`O�|6_l��goL���Zv�6�i>Z�]��]������3�q*@�'فN\���= �m��*�/��`~5�G�`�8p��g(�p!�y'�Ls�I;���l�
�?-u�woX'�s��Q��hLn�w@NHcY"J,C���w謂#:,�%&1�N�Fg���
1�ⳳW��yȚ)��e�#	Q	;�X*7~~�ԁ�߆R�мn&����W��4��j�вK�U��2+�����7j@ig�Ă�-g�����y���#���m�X��=/p9�F����Q�,�w����6�Xw��@~Jl���$r羨J��P ��K@&�zg�ߺ�iyY��2�X�i	I�<�Q��0o���:k̤��E��>��oYL�L�
}��޿*Ϻ�4Ò�w��JR�:�"�r�O���7�\�j5�ο��ŽMZ�-u.�7E֖����^+�V�,�|��/�I�s'�V�'���Ye�]x�w^a�|{�U�7�ڲ�>Km>X�K*���}J�W�k��"�0!/ )�,�����#F�{�J�n�[<���^ L���`H`Ȯ7hZֺ�)����]沰�I_._�a&�5,$T1�(<���M5o���
���M%%3��B����{�-����<����K���P9璍l0���1��ҝ��2�N� lH��tg���S�����$*��nHs��D�;�^�şkEwO�?M��	H̯�v��	�������
�20��9�t�	�μ�;�\�C�,`�h��uӧG�9+z�j����LMt��FIq�PC�r|A.�R�,��jS��^o�2�;�U�}��̺f�L����o�t*�L<��������1w����lY"�SI^�����(OT�ګ(�?I:
X"4�$T}rXz%�y��*�.�e��ED���P�'��ˆ
Ĳ2o�D��ʓD�k�E��Fq���a����5�h��B1T�u5up��"yO�h� �����\�?�N6k���wm��ZØ�'�1�HQnr$�\�*��ZZ�{s�9�@�~	L�.��n����A�1�g�x��d�e���A��|e�z`A�����$V��X�i��uV�a��e-|hS�/�F!���/��
+��[&���vdRw"l�C��6*��%��#~�u+
˶�ؠwx�����zK��4a̽��g��K.ڋc�+R1�2�s��{��ɔ��OD�v%	���u�讌�|5�:N�o��[TeK��¡K���_�xG�b�l�?0e����*Փ��nt�"N��E=�!YIhʌ:b/�i���)�	1���R�}<e��+d���v�B X���v�����U�^ڇ�}eiݏk ��T���<���y�Ah\š�1�ٔ����8W2C��y�d���;�z��²	l>����9��}5��15SJ�����_�7���d��X�W��Bk���p�۩	��k��"��^��f3�6��	:xHy%��=ya�J�/�����Z��2�z�k�r}03���2���m��+�#����r<\,G�{7���%��Z����������c����`�B�rD����Q"�C��QÝad�U�=��9Y
�@Z	�Mk��.b�[���7Cv�?Ϳ���e�K.G���(�vM�gnm��#@fAG�D%cB�����2�WQ,_y����Ur�d !�O)����c/�AjТ��^��c+5��cΩt�sD9�
ܾ0���`��ʧ�NSkL��QI��]��1[�;n	>R��s��i�r!S@ ��G/�O�OP�X6N{��l�u^�m�T�}&�?+���{^ŵT���r����L�#��5^�8��y�8�Tß,�t�ο���Ȅ a���}#�y�G��Z�b�����G���9(;`�) x��3؈�hIL���V�RE#��;޹RQ�g���L�;��h@���%�5,�\��[�NW�sa�Fb��u*ƽ�%B�O%��x�����'_8/��J������p\��w��7��o5;:��ZZ�m��� ɕp ��7P/4����یq8%��C��Y�k����U�@�Ӕ�N�3 �i�ñCe--EK8�?�/�k���C���Ήb�f�N��K�+P؆���}���J=#�'���[+ʝ�����i�D���Lb�6"�X�ұ��)�E��3)��	���W���Y����6mҶ3�i�	����~��=��P��]B9^t��A��ka��A�p�[γo�T�h�;�J ���q��!%UC=�:ԗ�#"�Q�)9ᰲM@iYH[�E�d�JG���?�$���sm�:�Y旟_z�	&���7�h��G��a|Z��1�_��h�H�e'�������:��i}�˒+$�A���5�g4��n��s��Â����'�����Hpw $1���\���?�IX{�����!R0�'�C����ʦ)�]�U�q���w�C��R�i)�9LQC�yr8����hq+��t|k�S~����lC�i:R��#JR��������J9`�!h��@o�.�tb��h�y�Z�Ɨ��1e�`�>�~�Չ��\[;c��w��R8t���l�"��5"E��ت=�QoS����Tx�ˣ�r9�m�B�v݈Z���� P�<�,r��;�T�;�������K#��l3��J�.�O��p�B �N�t�О�|��+��eC[_N��vJ s(�Я-X��P��q�����iv+ި#U���̐�'��K��G��=Z0�� sZ6���,=��!y�,Q�������r���i��� s� E��$N/iV�����;��-Y�&�f�e�D�ayK��k�^�0���D/�Z��UG��b�GW�Ί}*<�7I~��oB]���X����n��}��[�� BzD��ocC�@��J[�!A���n�����-!���9�>��匝�:2�����AU�����{��n'ytQ�VE���a����2��z�,'*��|����f�ku
�4�Z>��ܜ	��ͷ6a(J�lc��Q8�QVU����CS����%�34�Ǧ�z�K����\���?�>�*�ֵXU�F/�.����$CO���г��C��������_j
y�Xt��M�fiqt��׶����������~�\�'s���zlP-�ͬ��B��[u�WT��t�3R��ne�A���G��a7��\k�
�X��^4������_��h-��J�=&��׫�<u�{���#H$-�W�;1Ǌ>o4��A�s���`��Qs*&����м&�.�S��w}�30P�P&�t�ȂyrP������;ip,���݇�+���b�r�BT�%�Ǣ.��r���w�z�FT1�nߴ�Q)�J��;ʛ�K��;0PG�-�����^��|7����Y��訩�B�4�$�,�N�,c�Scb`/> 4�!�E��K�1�%�+�Hb@�{B-�- ��55ݩ��W�v��y�'��*�[t
��;D�� �ˈr����3�����#�����B.A7�-U�Ս6Ym<?�$A9 ���0'|�nvAu0�z���A�h�6���8"�^��U\]�͓<���]����|Y�װ�Z'��L�Ɔ�2�����e�Wu�ņ5L(?qƌ��b�}��᳣sɿ�T\9>/��h�y���O�-�n���}g��[�|���B�[�*�O�9p,)��/bgob����^ӧ�<
E�l������r �e1���� �S�^�]e��9�}��b9�)і��ַu����
�(�
�P��f/6�����w�$8�Y�iX��RÏ2ܷ�C����<AA�Jn���S�nYd'�`݆��9�~�co,�f�a�)㐗�ɗ��:�BV��:w�l��H�Ţ�.��$���=��j/��
ϲ��X��	��H�f��^Z�p#w4fd��]E��'��.U��Cl���D,A�4�U��m<��!�m����D��I'F~�V�Kk+�(�vi�ɼ��LFs����JH�f�=� �W1�{Kc�S�`��*�xfKP�x�Q_����`Z6��`�`���:�����!�^T11�@-�y_�l5w��nv�3~/8�>A�A��E��.SjAFvi˰*����d���ʛu{�� =�ڹ��bl�U��S`z�₅ �ӝ�G'��Ӥ��K�^�	���!�D0����{�he����=)E�Y&����b7���C{Jx�0�n	5)��Hq�(�uY�bL��o���0��[޶����ų��z��n��دn��Z4��he�8�`���QP���."R&)!	�.Ja*�=����@�gR�46���b~b�5ta���C*�T|�����,��;6�f�*�Kh��-B���U5% �����14[}	���]�|����49��Z+x�<�)�fzkY���n9���䵳��󇧙C���W5���c2�݃vC�ۈt�+�m9z���8����q��-fp�ͤ��G��~xr����ዡic�<o���.ʅZ�K�Eɯ�\0�?���Ft��<������&}�k���5(��!�A��+}6�෭ZQT-G�z<%��#��`Oݼ"kHB��ʁ��p�ᔅTe�g((ٵX;;��yȁS3�U�z�AD�v�POҌ�)����_���oI�c��uZ��'vyZ+K��C�Y<��A���"�2x,m��so6�������R�7�R,$�����I��4&.�
�|�+��`��T4bOM���h
%~��T3�v����󢀷�Kk��g���Q������H������^8�!$�������'��!�+*�I�Rl}�Ҝ!�M'FW��޴)��ݿ���@��3@`����Jng�NQ�	o�2��+?���f��s�sN��*�[�8�Y]}c�-JԞ5Y�E��L��/3BPLhRԴ��Y�M�|-���aGBC��J;!��B0-nu�^t��ĩZ�ٰ�T}�g�ƌ����.�Y���;�Uȅ��P�'���~���s8b)��8Х�6ߋt���'[#̛�ŀ�a�B�%�թE��b��G��]�.�Uk7v(>��xYl%`Ӥ�X!���zHλ.����h���fnJ�%�.i��AD�sh5鮹�E���?���s2�����JΏ���]
{_3M��?Ζth��u.�a�B�ϝ�|�V�/ओ�c�/�(9mI�/��.��Je�u �^r���o����ĳ{�1I�GBu�یȢ0ˁ��-,��*�q�}�]��	u���p�V7ږn�C�����5���㴔��"�WSeA�M�j�)����q�f3/��b�q��vK���p> Ц�r��8FAӅ|�Eē}02^��)aTAJji��&�=ߩ�>�����Mq�@/�dd�]���<sY؅`+o)����B�����6�
�
Vlg�8�R�=�d���M���2�I64�8M3M�۠�t�m��vs= _�vX���Յ*�8`H Gb��Bn�K,n_�^�ԛ�\��8���e��#�j��2�M^׺�B�q��A���1o�"�܆~���?UF���V^���#�d�����a*�M���*mW� #�w�A��F�Gp��%&��ԦG�|mJ�u��^�T���W�b}B
��?�W/��l���?@k�v➪��Mmc�Un�O�=o/���R8=�A�?	E?��u��	��d'�UQ-��X�ہ�ow\��ܭ=�adrn��YK
P4E��J:A��j/VW9����&�4�Z�H�����B��6]����g�Y�r[%�����]g�Y���L�}�0�}Xl���
T^���~k/~�{�߻%�8/ȧ��6Q6�¼Mc�&��7��0������CEKLٯ�q�<��l��0hX�J=RH߸���V��n:7��6� �b�w��>���¦g%�j�xY�I]ߛ
k1',�F_E�M�\�<�"P�h�**q��Jmt�G�+g�6V������f���߆�q��{�O��������=3q2���[dIȖ@y��I�A����58)��ӜJ�l��~A��Y�v*^K��[��n�<_BF�t��a���]�|��LD�y�L�]��3�d|��A�!���㰹-	����T��Zk����^���nM#:��l���=a��v�G{#ZEE�SW�~7���wz�E�w�#��w؂*��Q3�S/N�=3ub3���Ԗ�R� PL�j\��~Eda����`�\�[ށC���c��D[�k�S��,	�^:([�!fa���z'������A؀W��so۴h΋nŬ+�`�i_���`��-yB9������ⰸ���U\�}v$�0)N�2��t��E�������_�BD�U���`��v�J]�E���^�L�,�*ȓ���J"�gm�gӊ������ �6c����35b������	_;�`$�M\=z´r���R��/����׷C��jr�9o��4��:Dv��Ilݻ�������,K�2�* ��vXS�a�������FX���WW�ۄ�r��Lq`j-�3��<,��u_�n|��I�p�>U��K|{���
 ZRV�0�܎����pe���ߍ)ȅ��Pk����ܱ����)��TCf��dC)�v|��Nn:�����U�I�R��t�`6�����;!?C��߼dl���9=����ɻ�X7������菒�R�O��Z^��A�C8~���	g���Kv/�6��fՆ>��Eچc��ðU���Z�d�Mu�\Y�?��;����#�i]�W<�@#gCΗW��B�En�jA���ѮV\�3'�r�zC��vx��[Z�6�+�@G"0�)�>��y#v g8JL�~��Q��zF?�ұ��,����H��0	�2�к�.�D�!"o�g�K��b=���׷�����œ⒚_��k�n��G>�;u��x��Iox��3C���O��l��g�Y��qcAIS�:�$"���o�%>b� C@bkq�5L�|���e�<�9���~�Q������CQ����RZ`��j�T;
�dO���,��H$�B�)�xecgd�h6]߫��V�I��ϪU�i�Y)n|��"��B��ݕ�Yb����[������Oe�������Uc�B��,�Ԣ�S���V����g�&u�K X^�a��Lr�M>5���(FAI�JqC�1�Q�ֈ%���E띓y�9V��T�%��̽�/�`!����L{+��cI~�"J��]V���,奚m���k��OKG�PU�*�.��Vѐ�lh�A.&S$�;�V��!��.w���\:ݸ#�{�EŌ�q�l���=����Q�*Y�~�����ə�^��a�e��jx���[�ymXx���q!���fs�V Z���#9�C�3��
}ʇ���7�A`\ԝ�c������ٵ"B^��e�v)�W](����Ί�ߔ�Æ������v�%J�&�Va��Z�V�#�(��C�5yU&�}r�v$�gχMy��r)�/-���� �<�	�&�����0�-��L��=��{���#�N]�	�.�5A��ԧ��#2C�tA�c}�`����$ 譩���Sɨ�$n��:�FVy�^�S�(|�����R"8I�MA�O��6@�󥄼�/;��g'A�E�k��	��_n�6)�޳)�B���,�<����w3r���B�+e��/��a��K�%���a�a�����t�֫���N�'�09���Upɫ"��]s��6f��d�j3�x��*�����Q���Օ+#�<��6��=/��B�E��e���C���E�ճ��e3�&vN�~A��91�qS�GbZ��j�4[��B�?.9OH�@�1��xJ�r Z�4�g������T8<be[ڌ�犽���a�ُ:6��8�w�Y=�>/�:ֶ�)�Y�;��n���~��s�VzYQ���>]�2|�U922h 5Kޣw@4�fV���7����e%ʪX���v�3 z,����#�n5L�,��w���YQ(��n�=�u9��
�E}�D��l3>���͹k��Y<�����>�d!��!C���}��+��]�Fk�t��I'�F�w�>��\ϣ�PP��b^�ZW��MN����r�\��MI���x(���:���_�b����lv������)�1uI�Jʦ�>��Co�b�x��P���kAb|p��S� J�k",H�ov�x�S�
�B�ɞ^mn�}s��8�:ݒr"������x�! �Qy3�Y/�?��;���g?X��O8Q��:�Z*��dp������lg*��@�w_�f�Q��x�W�G]i7o(Wq���Ͼ�cSʁ��@#�D�7��z�j{v<��7� oBk�J���Tw�� +�¼�0�-z= �F_	���<Ӝ�-���F&P0��i\^���e��8
H����\�?��mz�@��ۢE�b�ܒUlrf���`�)H��Lz]E�*>$^))R��N�gޡ�ZE�3��=�<�i�,�:�U���i�w|�H��Yf�&��S�Z	�*�~�U��4��A.Nu�d�Bc��퓽[�e���� �A�%4�����~~ywF�8$�	�P:�dDLQ�o��D=a#��\8��#XM��-��R��4,s(�����F��6��?N"4���42�H�0�{{�G.��o���X�VbsO��;O��E%�#\h�N�4S�~T���p���9�V�~����/�Kt*�|dh��eF�����H�5k���f1��|
9�8)%;(C�s������	�<W44�wO{����t�=6��<�Q1|�'����-P;$�J}��粙	F;6 TC�#���i���i>1�z�mP������W��MXy0`�� 	ڱ,%h��y",�>P|F��!R����J$wB��w�x�aB�n.(��#����R�WU���Π��j5�Հ ��"6x�����sb�D�p=�$u�?��������� �n�Y���O��B�U��g�;�P3o}(`^���/�ɰK���U6�N\X�jՌ�s��R$X� x�&��3�_a�&�M�$҇��78k�}NÑ'Q��(�R��uBl��Vz��,�)���咛����������2E �w�̉Z�D6Ӧ7���X��ɤ�/�����A��Iu�c�~����1�5f;���{B�F�E�����#F7a۵��P��,vf�,U�Uz��	���ν��s��MX܍��
��a4���x��k	O��*�2���i�l}yy0j��a��)��x�*�~fi��\B(�B�ٷ��7s�����S^�GϹ�Hp���п8��ϵ]e�?�B,�v���&rF8��U��,N�>�G�9�\汥O�G��k�{0)��U&V��G���O��O[gxD�L��+��y��v�=�K0�z�HQ`�)N��h]m�H ��*�n����� �[!�svnqK��� �#�xB�أZ[����_��G�YͲ�R�/77�Ǻ+�<���KX��������OT�(l�9=��rf	��C�帴���;1B�ճ�����9���b/��1ą8�>A��3[�uF�[L�x�#̠�����%#�����|��1DC}N.�� ��$Vi�[������N�O����Bi�4FD0����@�x�$Xf2�GQ�{�oi��g��q|3Ϙ�?#Ez1O��}��}���r��Ҏ٫��t<<����� ��a�`����<�V{��L��]� ���ڍ	O�y�=���WLQ��ocYx�L��b �.j����E��z4��+")h*Կ>�Ct���"��`cC~�oA����1/�=@�)~��~�A��S1�*��&�0v��k�����>ߢӐ�G�[{��>�)���<pP��a����G�*9'�c�h�d1ct,ZoO���o0�S�ء��{F��?TT��#,w#, g���8��>��}*�mm��-���6�n��
.�^��->+5�ߟ\��%�0磝 u�t�<��/"?�8�abhC{����ɝ<8� .=.�}ExB�'��k��r�%��t1��&�zK��X%+�1�i8�\�?����� �l�OG^�Qi4/�h��N���Fk�z4<��Z	�ᔵ��?��s�v��< N��~��g�н�"0�"����2��vܢ��r��:�Ŵ!D~=�=D���@2��jZQ8�CS-�T��{]-%�(��@J'�F�%�!�t.�����:
C>�y�]�T�9JL�0�sC�����*tB"�9?��|/�H�R�M0�S��w�܈d�+��kUg j�e֞�jI��7����G�ErT��>��
D���_����/XRի�S�.�+��߰5G�|�"M/t
bk}����y �l�M��'�ȳYq��faMN�� �T�l�e��Z.�r���662�O�ZD�n*HtG.N�;�,Yߙ�p.t��-Ҽ/����+���-�R;��#Ma�����%���aäO��P�l7׼�P�V���߆�	�'�M�]� �"O�}	53��<�B;�c�jY1h��+��ǉi>��ɲ]�D��P�:|�?�v&6��+).�V���p�9͠\�^���DZ��O��Py���� ��9���Ey��;��zeX������M�sSx��X	q4�bD i��=%˷��f��� ��ǽT�g=06��m&�:e���;GH����2���k3���~�\Y̚ۆ֊�9#���˒�RT"��%���R�V���A�ر�35n���[Ԋ����dU��!�WTA^�H�.�(-Yp��jAk�`����c
p��w_�"q�4��/�kK�3�ҙ	��6���Q�&J2�/E:��e@GW0�����Rѭ�Lx���`�b2�uRB1zP�Z�k��-�)^0`�y�b��������yȴ��0�\	��=l9c�Q8�8Q6���D��{;	�$Z���Ĳ�z<����$ܔxM�>8��@A��R$�q8����-���¬�����e�N��!y�ܯgF3�_�Kt��a*TkL��G�Yj�D]��>&^��FF�.��N���{d�}��i|Y�&yy>��t��oWR�V��9�mMy��fL-0<Fn�{p�J�ZZ���BC3���=�\p�)�v��Y��9�b����zsC鳇XX����$��h�:x0D+���fTZ_�lbP����P��YJ�[�T��B�֖��,�^�_m����e���2ψ@��؛�Nf`@$����~a:��w[��ׄ�B�ܕ�S�i��VW	�9p��>�Ft9�C(�#aMCF�;;5�_�M"W2�h�N����(�uHy=V����3���NS��x!�����6��� ��W%c����ƚ%���*PZ�J�CROR/eF-O]�ޅ��27�l@=�&���{&����?Z�
���9.�E垫'{�(ŉ������.ӻO�j���\�aAD߳[�Jǂf�]SjfZ-Dj
�C�)�N������Q���J�#��}E�2^��0�~�% �?hw­8�8Di��H!�!�~fx���r���M2,�tQ95+0�	���-�P���2���vJ��*9����B�b���c�ݴ����m9�2����7C�CgF:�vS��,Z��OU гמ7�٨�m��`9��Ev�zϛ�a����}>ԡ�;uʍ(��`�
�|%�U�rZ���JŤ�?�`�B�;^�zUd���ʹvX�Z��c�:(�#�F��FFG�O�)�B8up�������^����G6�C�\�ٔ�4b���5"����{��Sq�~$�Yl��&�¿��_UIhJ�*D�8:oȱ;c��~��z+x��\;T>cL�a���Ug`S��@�^�}y�x�.H�D����--Dh�� ��N��)`�_Ay@�U���uz���;fy�4�+���ֵԹ]_���5���@)Ҳ�O������xp���R�6$��r-k�5��leV�J!����&WSd�
-�&;s��{�c���_��s?�j߲�r;M�xISG���i̬�L�(�xvY�J���f������@�{\5n/B�4 14��6�}/ũ�0��wd��E�N��M��R9П�9�_�q���G��&���fA)<ǰJ��QA[c��T��}B8{�lH&]�����("@�`�����l| ��^&u\�G�^��� 7mBM��&0�g�ND'�q�Z@�����A�6��n�Օ�u�Y��N���#��>�8��X�GǈJ36�?���ۤ��YAQ^�/��G՟��-KL�hcIjNǪ��"�;�;W� ��F���H#'#6�I���%����q��/ɒK�K��5��鞓P�39v��Ol��*��	yو�V�lf{\��ȍ��{�Z���2��������P~c��Kr+\�QM�fa�V�蒠J�뫲��r̓������_f_1<L�?�q��EO��l��,ʗ��42õ�Rl���O���:���3u�Clg+o��U����1�����3����bG?�%k���e$ e��/5�\�u���0+~�>>c�i�Caot� ��/RO�I��0��\��ߴVrU4��b�>��lY�;a��m�ں6$���Ft�:`WR5�/����͖������M�Wrb�@H��sD�RI4s$ߞEZNQ��s���ܸ��h�=�I��ڰ:	Z���
�ƪG�o|lnŢ�[�Հ��S��w|�|�b�
9�'�V�<�ć�ᓕ\������^ �
���Bl����[}n8O<Q�E�U���`�|��_@�?��;�Q���W]�Ý�'U-1�K�I4�H`��Ϋ1W��~��^Κ��ძ����ު�As����W:_�E+K�,�x89�/}|�>��ӔΉ <��Q#l��s���Y(1�=KiX�'\�_�v�
��DY�JW��O�¯r<�~f�3yG���6ƈG M^�����4OH�D��?��W��u�"X���.T��IIH��<S� �:����G�x��?�?����y] 1�-��-�UT�[ڬ��^!���%GK1�W�֬�.�H��|G��}��3n��C#�AC
pF��.]�}S� �_��b��:�&U�cQ�g�cTu��7?u�Q�@�9���Ă�Z�67S��;�q���~Z��_�ɋPl��w� �
zl�o��lj��H�Ҝ���D����o0s�t��a���IC�l��h�:t����,�J���yP� @b�Dݎ�u�_�F�ZH-X������@�w{���q2|�j�4`�ab��6}y���#wL8.B���("��U�L���Y�;H"ߩ�d�r��z_���
Q�M�y)��[��}u��9���G4e���!C5�5u6���]G��)̔�Gc7!<�i6̱X�CF���׈
�#�ngy.?����ѿ�,��m�c�Xτi��	�Q�R���c����犉`��N(S�b�i1~���W9�A�}ӷ��<�Y�D�6��z@*ɏ'H!�Q1��a@IDt��"W����6މ���Ӭ,�L>h�	�V����T��~�� ר��C�p�H�O���������E�W|y_P׎��ެ啢��T}�.?E�%֚<Ӈ���O�%h�fg�1;K�>�	���@K��o{Z ���B�XT�?���
�j�ƻ�!��l��t~`����8�~B�᦬�8���i�?�E�5�ܶ_������W0�~�x6Z�k��g�]��?����u��6:x�Ү�R���y)� p�BKЊ�(�(����9�@��$�!�<�����'�'a+n2y���BS�� (lf����I-���o����U텅���x�V���u:T�ZH�Y:����Q��Ģs�iCO�0�F}�q}�Q/���i,0�F��$����l�S�ml-{Y�N&�&R@�J�%�;3�<�5A��j,�Dc�aS�O]����?� ��CZK��-L������Z��?���P*l�c�*�jY&Kl[|�gdS�am_[;10���]�BN��n�ņk"���<� ON�"���W1��+����N���'�#�$�cC�:][��P-^�R��9m��<�=6vyX �T�Ua97�B�v8a�t�x���IO2��gC_���A���0�8e��1�P���s~�.�`J�@+8k�[U�4!uB�'D�� ����g1��"BZ򻒾���I�O��,.�_ �����M���*�������K��f�B;����I^��?�f�M��UM��6���4���V��m������;ޝ�d�o�[y~����һ��Dr��T�\ov����-��ֻv&mc��k��OE��Q�
�'�� :?��ց�z`�j��� z ��席�1)��]Χ4�2�,4ԉ*���ZzӬ�������SV��-W�d��$�"��t��8݁Vd�Ek��.�@9o)���z6^\�`�0��C�����Gw_	:��[�q���Ӡⶸ�;�Й6Ihfa��$��{��6��c;��>Ytc.�m����m�:�I�������뱠�#��!����jF���+�)D+���RX.+A7ƣ�T�hϷ���(!�,�s�{u	+y1�~a�$Bs�gT=h6HRSP���'=��B��E�*O�=XU��\M� `\D@ �S)-h��U�:��{���uL4�9�%dn��O�^�5k�f]�V ��|If����;q�������B{�G_�y��`��[�F�+~� 72�D�s�5����V6>�H0��<U���'t�=� �	M����ګ�&�0 �e8~����MXy�BNi�-�}|�̒�o�6:�c���_��e\	O�(���"����E�~�����jL��x�D�I��*;@��!BbviZA�<	UhO˧ӻ6�h����*~�P�6m�M`����p�/�3פ��W�v�(P���UhM���p�)��e+XQ��x�x��1��1��|j����s;���?X[���[�����^[�ηԯOL��[�Y�!������M�B�3ȁ�N�k"2������79�g6��2������@��jek'O��v���y(�v�~0���	�C�S;���[R�k5LQ8*Е=��(SY�Y�m7���D�]U2e�LӂW �������ȥ� �Mѿ�R�b��E	�됙�*((����������e�5��Pr|l�����2r�^�o{�2��ɉ�!����˶���y�w�R�E.1�-.۲=���?7}�P��Jy�H��Aq�%��{E�cx�����	��.�
ZF���I���N�S��Է ɜ'��W�k���C�K6E1��UG���CM�_BjXQ�Q��0<�:�F���Y�C��7$����:����:��ʰ�^Q�~��+q.W�����}/΂��}Rw#Q[Ie�X埀���p�n_�aPc��T�o�(�/m7������,�G�Vo�?�ﰿ,��WP�zK����g�Nݶ��TȡQ+X�n_�؍�(�a��ʪQ���n
y���8u�;��<�%J� �?�k�~:Ғf
�*:Y���;%R�)bu��dBa��uV(�Y��#�x�ˋ&���#����jn,���3���'>P��L�ȗ]b�A-����=H�N��R��u�� ���´u���h�w�NF!�?!�~oP�͙q��_�k���v(�|��w�)�ò������R�q�<�.#Eȼ�N'���2.b���`�i���yzf�&|�8(����7�u	P�M��f�go�0>��\}�Ex'�=��ʃ�u$���~j�ff�X��N�m�������ܐ���&�e;8�>��.:Ģ�˱--t)K������=v~@!xG�����HINDm����&�'��o9vԡZKV�`��J�Ҏ!E�8�k����I�	��xuxbf$T�Ġ��x;"�hM仙�����v,�=#D���	���t��4������T��.��5�5s�J
��8L#�$/s�s�p(_i3�&h���sE�v�[���P\+;c�Y�Y@}��߿�d��.w�걻.wrrr	���Ҍ^؄���De̎z�����74_^%�{f�9ؖ���x�z�f
JL�)�@���H�D6�N���V���\L���5���a��|)���c5�c �2$�@H6�LT�4TW���t��>�i�����T�4�R�#�;����nm��t�����U����3����s����R|�4��p�^��h��P���1Ê�4R:ҡ���r8RW��q��d�����f�;�=B����q�p{��4N�|qbn�d=H���}9�ۼ��1M+��,�	m��m������M5jl���Z��`�b�Qa���A;�iLnE����js)֘Q�`>���3��Z����uvW��;m��	L�Z��쉺=t�w^�s��!�U�Z���[^�|��,9Y���'�G�
���F�k���,�ټ�^OB���sjb��ԭ���Gv}�Z[vy����a�>���l��;Yi£!*ׄ!f���$|��h3���H�wN��V?�DR#�|��4�Y �j��(�Qp�Y���v������A��q���/=��&wG7WP�uz�SY2�{'��(}	=��(tsؖ{��5���贳6R��T��+�Ow3�B���!Z��G��7#�kF�X�6�+t �>�{���jŘ�+m�p=.�_8�%���-�͐�?i/]��@Q���7��0��1������i��SfpB�(����Y�|�Sb�5�e�Q9F�洞{b��+�Ќ(�m�yÆ���w��⸳�6l�@{ؿ牔g�"B��R�';�и�u�I`�Ⱦ��JP�P"l��-�A��Z!I�ZHC�ȯ}��]�j}.q�������d;�4T�nK7�_��+��.�4�V�Jʲ`nfi��L���H3��_�u��}�c����[1HȬ��vM �T�N�$]��Uݧ�-��ʙ��4.Í348�m�[˅$�l��$�r���~�G[W��j���f��P���/���t9O���f��->���CBH9"����*�m#�L�M�^�gD6��/�n�'ȫ�X m�{��?t��>-����}�'q,���~�1d2S�"v�ܶ�,�ۮL��-t��D�q����u:g��Е@A�̤�p�W(�/�ٿ'ŎV��Sl�T��.:u*�qU��[jvP����p���)�.����r����P��=7�𮤱7T)Ɵ�=k����D�hP�}�ZO?�1\{Ӳ��v�W�󜀂]%�P��~���<dx��|U%K&٦B�?!S`|�=$���!1��
�W'H(��Ow����]�� ZGD���`'�b��X�����YZ�o�ա��Hڭ"�~O=�YM�8���9h"�N�����9Г�^Y�l���ݺ��@3B�Ɣ�r�8rhݵ��� �ˉc�a1�y_�e�	�H�鐰=�����f?e�W6�>5+�յ��tw��-���v�V��+�_��!�Ž$M��6A]B�(n��~/��V%���F����L�QO�]\��tS�V͢�`���F��x4T㈖s��҇'���b��Kg֦��A�Nv�_��
�ee:����ɺŨfa��K����'זLRх@T��~�=e�GEicC˜�)�k��E���w�GL݆�(��	�2�����.R@�i��	�J�i����|
9p3b�mmyI��F���}!q����GB��9P��}�p��B���?�$�B`̱�g̷pt��͝/|>�U�ڣ`oI�z����c�{}��B5N��Y�r�����P���+�i���.���t]h=�<�𒆀��IO�ҦY?�p4<����M�)��y��F�_\�@�P�����m��U���|!=���Ȼl�Ji�t,Ќ�t�XȐ�Wѷ��� �M��؇�����I߀N5�g��%��C4��/��鞱N*�:����f ���B���j�JN9�8��^��*����X"A����k���Ui�$2�o��?S̽Mu1�t��N�e�g?z���k�U�秇R��|��u�a� �!���B�'���#čU�a�������F}���
k�G���/U��Wi�nF���p�'������ ����G�\Z�u>���3�%�֧%sr58_&�G]#��~,;<v��٥�k��~�9�qSF�����{�8[�j�	:ʧf�V��ְ�3L�9��GmC.c7��L>0�8�.�H'y���v$pBK�J�P��IՓ��D�fY*���r��)[ٹs���
�U�h�M��r�:��@{�,�����Ϛ����6�l�[�9rHo�i7�<�k��eiL���1�E'�X�H��uU�w ��rޝ�H��2e4>+�����Ǽ�r��9?r ;�����Ɛ��b%b�U)W����Bc��m,��5h0㛟�67�J�?����nE�m���?ӕ�G�}�/�HXêE�Q��Ql��bB�d���+cҫ(�Xt3,[�AC����R"�T����	�ѤNa�`�ɴ�q'vB����+�-@KD 9����ﮊ�RׅvQZ�>���W|K;	��3K�0M����m�GXԡ����e]��e�
jh7�L�����xw��݅!b#��_��?sB�Wc��7����s	�M!��Ћ��)6�P����w3	Xm�[q��p뤒�,�k�4��od�"�q�bm�'�y�4�e���!#N�*�"� ���sT�Xvb7w�+Z�X�_�&��K!��lƟ�q�t߷V]G�4i6�U�4,�]�g1�b��E��aiڅ\o��o22��K�����"����Y� ������)/
[7;�2	��q,`�C9M��6]RT/�x��˞K)V��h
B*�A�B�b׬������H�����g�V@A�yE�l���Iln���,�/g	ťP�8�ov��P1~�@ð� n7�ם_y�X����,��Bɲ�7�_Juԥ9��&"(��7�� �������q��&x_wn�C��x�1��&�f*��i�ц^jF��6w�24HC��q���� �ȭ�S~�\��t<���iF��d��/�p��;��0J>ٕ�Z��S��8W�YQ���Y�Qxe�0KcA�H�]Zf2��ڢ�!����j�@ת��������
���6��E':+9Q�v�I�H:?��4���ۇ<$��ѐ�2J���.}��n����,�5
���Ql���D�وT*
Q�ӈ��J4���6�f�3$%��Ȍ�o�[�
�2�W��Sz�p�w��}�����}B��$���sdJ�����/��s���9�dQ�cH��~���M�Cs���hV�K��؄�:�v�a�9�������h�9a-s��g�*=_���*�XIP����V�2���M�ӳ��rR�3h|�8vN�'#o���z` �Ԣ(}� �&S�l�dntO�iƗ� t�W�'}u��Q�G�k �C��;�E��A�ȏ�&z<�|zwTD�~��UO�I��q��T�f�t,G[����j� �dY��M;gAb6d'J��o>��B��*����� ������J秪��YI���m�o���Rt-}Ci햍���|9�H��o��jm���?Ƌ{�!AR�^��0�r����؋�g��?p�uS۾}�� �!Fݐ����k�� �S��iq�����>z��1k�lJC�C�<����BPg�&��)��Z����[�1�x�#1���Jj����j��ùJK E��Zt�
��-+	����Q�ЇXi��w�) .ˌ��l-�T�;&A8�51W�}�	�5��ߞO7�e�+^͏b���LU �|�^q�L����n?1�l�v�Q���w��[�i���IyO1V��B`�n˨fp��Zt�M��Y���!��o��D`����M�hk��`���e��L�r=ip�[�
,���c�Q`t�{0����) +4��?a P��ٓ�$DIc=H����U�I�?؁X\%��r\@�2�j�4����dB�JlG����9�+r=�i:M&�a{@��7F{��)i+V\gI��@^ǫW���mc`�a�������w6���$�. ��R�q����F��V�%�7<�81y^�Hٞ�����R>��w:3>k�q�4�f{��X���v���B@�ϗd�N ��+�H���:߶��4bo�LDx�>�Ĉ��oB ���6�L�1ISS}u݉u���;�Q�����@M��X� ����� )�k���qb�.�@�L�B���vK���+2j�<��>��$񋖀v�~���J�F�j�����+�O�=U��E
 O����>�/P��%<�{~�:�ú�\�.B�>:���N^��&�#��0��^H�D� ��p�Fi���uk�fIߑ���F�]lt��Ǣ�1o²��ﷇ�da�R�ZӏL�[���q׳� 8y'�u���p��2n�˾@������������sK#�'[&�e��Eq40l�Ҍ�	�\42�OH����U@�e#���N�v'-	, G�̈́`^��)+�N��k��Px��`�d*����N�2d.�4<�)�pfK'�,v~�ҍ�������6�)}y-_�z��Ƕ�VѶ=��ğ����@+ZA&�\9VO� ���F���r@i���΋�$����O���`�iA�!��0#�ތ�O���P/:'���uwY�_/����o��ƞ��@s����i��M�70����6��_�ڿo�#7��6���-�>�Z����S~$Mʔ;����1.R���0#�;�m3i;}sUx�u[��X�$$ kY����������X���Z'��ehns�����Vs���̌�-?�E�p��2�nE����PcTcn�F�;Oխ9b����f(�7$`���j�x�X�	��o3D��II?|�z*�*��,e=!�frG��_3s�&�/�#Ǝ�������
�� 8:(�Oͅ�q�4?�<)󧘁��S��I�6�<=��p}�`���5ݬo���y�L�ӭ:�k�� G���r<"i�MXw'3j����r�`�C��_��N?��-�R��=��R�_��v���L���+� ��8���f�Y��O�\�t�.�,��� �R���Vj>"�0��5bs͍\OZi�O]��b�!s��Iӷѽ����7t��m�ߵ|8*Z���</�Tls4Zl��eȞ͈l�K"{��(��n\�4��//�!�>P}�$����`���	�Puh�^�k�7�0�0>f���p�=T���;Ɯ^\|)i?23��b�yQ� �����@e$��U�F.�������"up��.:��������i�r��W�ɵ@���B��;���r4�04�x�-x���O恫Ʀ^uI�<@�Xcz�F��|`��h��)}�JٞY�����f�FTM�S���:��C�N.�Xa��� �*�������v�ϵ���}����:kO�<ݮ8��2C�C�*���lWL�j$-��Q�)B�^<������d)c�Ђmu�j��i�m�׍�b8���Xi*˩t@��e���T����"�IɃR[�/�E��v�<��	K�ا�s�����J��B�ř��B�=�j]���h}��D�`Q���$�G��J��0��RqC�XwXU_�f���0����5'��C��=M�	�Z_��k�ts�§�N����_T�<E9�&	s���n/��"��qAW_ʚ�)��0_L��i~a���� �.��5^��L���	S-k+�E�EЄ%���k��pޯLz�0~��T�)�L6���:#M�l���m��= ��n�9�L�fM5��?���60'/��`!�a�?�w�lV���~� ���(s�5=P@���) "�����U��Rw�ؼ�n˚���ʋ�v��
���I2�N!��������-&<ѺE6���Ѳ`��q����q����,o'�ȧ�����T�|�M_�E��M�v�ՎXgZ��k�� �{��#��D�bJ��m�8$���C�G��B��a5������S��8����5���T;}��Ƽ�!ѓ��T��!v4����ү7��}fR��Z����4����e}*]��yC{��]k�����UX�Pr3.�;{��|������A&L����[�����u@�2?����U*��s`2���t����/�M�U�2'٢�f�m���WK�+�zL�E�����X�Z��2�`y���8;��t��RZ�����*w��}�+��Ƃ�*�c�� YƵ2�aך>�`,ݝ���F�D�
�Y6��5��#�3��ϧq��ᵁ�?UץZoUM��,����y�Τ}[����u��j��s�5�'��Rٟ��.�û��p��(WY�F�>__�S�O؂��AS+^M1Ltx��6�*Hg=(b+����~���m�}Ll�v�v<;R�@Z�,M����	���\ow
�!�u���T��_+&" m�q�Ǟ��l����
o�n�N{�+��\zZ3��ʟ`ڇ��b��yC��m�)tV�'��<e8[�|�K5�IK�AHS��J����>u�ї)���E�Enw��7�9���4����&�j�M~FO�>^�;��^�I�;�H~|�@���K,�	��u��,(9q:�(�=�e�݉�{F~�߮5Uz=��;�)�L�,���5})�ǂcg��:B���Ʃ21�k��û�)�.�â���)���Ї��`��&r+��,���t���}�E�
�߅Р%������#;[JY�$)��+�z��1���]K�f>U�No��	�%��^��P>�
��L^9�Gh�~16���3����V�r�NN��ySZ[Z�M���>��_nIХpD����q`�݉]�$�/͒��L}�Ya� ���`/����]H�X����ܑ�c~�<�GI�9�xņz�k�;,M�6`�umꮨ����{h�N�d);��ì�i`p dE�r���\�t�{�;<Ir��Z��%Ȇ��C�!���Kꖹe\N��KU��x��3�Ql�l��v�t�-m����^����)�Q�C���	�
t���&o������^M�+oCN�n�q'��$:���~z�A6G�w2�\pt*(�}���v�-T�`ֿ}='��>�/;�J;�,����^^�\��R'�5��� �t��3�-�$�I�FXm���)���>����7�<����d�x<�����X�Y}7���BnڞS�Ug�n��<�G
�6�墳0�B��{��+���wm�+O�������r�������d��+���ȁ�A���}D��Q��g*��Ͷ<��s ��DKW?�W����"�R^�jX҂3��ĉ���t�)�H�B��&gΡ�sm��Q��Z1���4T��$�����<�J�������e�fl�(w[u�.��S��|�y�Qt�p��jd�Xg�N:��9@� t�.�9 9��v�R�j��>���+�1�詷������3��A��z�@Ŕ�\���Ἦx1��3�̎)dr�ZKO�����K:�|7��jtQ�~��Ȱ��-�1O�Gm�@h��̸�qZa�dZ�����W���(1�U׳?��f�z�D����P�=�X�(i���E/mz�}�W�|6��5�Mŏ�(l X[V2gW��P��2���&�a�ߓ�a��Gb�n��y��i��
wS>�f���Yk5<vR�*>���nG(��iؓ�A�z�e$w�s�i;���S��b��bm>�S������#	^��;Ob�Q�l@�]*3k���+��YmO]:�m
���{#rq������vJ^�ܻ��]ѕ`d&u���H�U�գ�8�đ�q���$���Ā��.m �޴"���SHD˺�Ix�P�/���3�v�� �4����#R��ޝlս��/��2ݤ��fӕ�N�.;:�Gs�� 9�騆���6���k[��By�,6k�d��hzx�:Z�b/z3M�Ѻ8��ݔe�x*�?TH(�w�M��2[ơZ�3���=4CX�o��aW/�n ��6�i���
��q��D=��T�!�N+��<~�0"j�* �(���Vͼ�4�
.Z�[�w�������d�D�G\�(��#/qDa&��Ft\��b׀��x@�(�aصw��P��h����dT�����Q�#�K|<o0����ǹ�"�Jy�=0�c0��Q�d������C����R��8�q	QUO.��+D��#ĳTK��!ۚ����uֿ�+�w}� �:)"�X�c����_@�2�ˣH���G�-+�V�R�63l/�pVg5ᬷ��+�!�>���*�7e��jG����nF�:U���䢏0QA*4}��C�t�����]�`~�6>B7"������jPO��b%:`��5�?�J��f�J���N/�H�� n���Gޘ9�q�-js#O�i껀�XB>{#��;l��c�u[����5��M_5E�`��0��~��Y�f����C�1�:�Es�m�fA\xtj;�oŴ��WQ�d��؆#u�KW�to� ��z�%F���1.a�+��~�:�ŗ�mڸګ_�K*P��FH�I�D>3�Pv�^B�B@�D�-\3��:[&�_��Bx ���_k!�m��u�������tZ���Y�"�U�ߏ9 g�x�7�j�&Ȏ��HcKf�,w��z���w���C��Z��Ei���܀|P�@�p��=����(i]���c�����-�)��#O����K4�����o���0���+����.E�,��W}�}��m�Z6���hSF�Knӯ��{"��AnBph���?�C9�cee�����⼰5�thk2�(�G��a��V3;���B�FJm��h$'��?]�1Ti��0� Ҕ�#�&<l3z*���.+P�u��#u�(�M!��	Ν?��e����� T��؊��S���4僀�W�?V�EM���~�;��	#U ���z��LF�~_̲3�4�<��RCX"Dd����K���1����>*����W��
����]��W��$� Kodu{��Lb�����@���t�����W�:|���mc�tN<w�TB��U&���G�o���[~��,6�I.���uƈ2��>S��f��u]���k��?ax�*�]A�gfU�iP����֜����c����ެRs��P�i_�sE�_c�co������&r���n 1�)�NA��;�ౚt>Y���߷)�[c�7�l�k�3mL�b�������e�1INZ/���a&ߋ����כ(�P��ᮾ�ƏA>	,�ވɶL��D�� b]jO>Sa�v��V�����U�Uʝز�-��c"W�g��N]�ݥ�/yz���h�4��\��N�f�Cj?�&������T@!�D_VJT�.�9`y��ץt�k����:�m�	O��@n�4�%��@������M�^�W��L���t<��`�:q�j)]�֘�`�
��I����B�X���[`a΅UzJbպvY��P#���ֶr-e�
���8�_3�Tv�3T����2�8�25�1�*�嬎�V�^�*P�J�6�Y��7��V�~KƧr� �<Rs��Ǹ����b�~Τ$+R:r�Tt�Ii���4�c���@�L�rT��54�,ʶ,4�ť�9[p��"�b�R��M^��)�3I�����&y"�6iՃԉ�q������D��Cjo�:�l����#$�%a`�eXtW0�Ы{����q^��[�k`� <y���$�j!�c��K@X��Y"�'��1,�Pr?bPv`|�����#����4��d1(���Hf	U
t7�!2�L��
��O�kHt]k��0�(�GV$��B �/ )E��y��Ayh�K��&�?���"8�|tġ���C.��V27t��%���խ^r���Y�.���R$�i:R���Y�� ��?}R��
	=Ϥ��C�E�^�Tpk�j��b+u��K�HQ��1*g��LvN�Ώ�0HK��z1O\���(���_�9ᰙH�RfWV����z
���W<~/�J)��O���iU�h��ߴ����{n7{�t���bmTۉ�cp�*D��k���^���VTHs׼W�}}�Z��E �7��W7A���}*	���m����M�ϣ[�˂��M&G�4K'I���:�R�-�`B��ƪ��	J����h+ۡ������Є�QQ��u�2�*ƛp[���#��a8�����^.��9.����9+r���,�M�&U7�ݬ�6XE뉜A��f�ؼR|��Q���{���M�D?�U�)oh�m��7�e�q=B�5D�ml��&A�����5]&U^��#�"�.����W�px��[梋�P�p�z"�'-� �B����d����ҋ4�P+\��^����w��+����t��	h���u����c)+��jEk���HD�e&)d�L�2QkJ�PR��s��v��u/�?�,�qhl-2�8�
���$�&L�T8�?�SV�f���B��f�3V���ۛ�Ci�[��
oE]->�#��eǗ*��pl&Ur��� ��Hv�l�Bn�&Ė��F7�܌�r�V����e�R�1cb�����¯	ik��u�dƋ�/���0Rl�84���{��i����E;'�<��J�bZa��+���ըtx�ru��,e�˺jN:����5ٻ.^�W`�e�ˆ2w�F�dJ� ��
�Q(%"�T�9�Վ4G��W覕�x2EB+}}Q�١���ss�>�vpÁ�/Dw�c���M��w�@H�D�kfk�=�����=�*ˁ�r^��o@.#_��t�I�.9����(7*�ݘ�!��Q�Ǘ��oy�'��3�,8�}��R����Ky�s�,�g�D\1hKG&�M������c�Фd��*�NU�u�sJ�!�n�3���=yl��vn|hǭ����ʏeN|ۯAt>ii��q���~��!M~���I^��9T0�ꠋB�@|Xm�W�I��Ujaub���N=\ecaE� sM�z�J$���k��ۘ�)��2���E�l{�[5��S���q�3��j��VIL�����s���o ���T��VE�۩�R�Ж�OuV�1��r,֐�� $�[�Eff$	�>`����I��Һtn
�������Ԏ~�n��!�yS������ߕ%`���~���'���\�A��������V�N���ת�ik���o����������ayݝ��?����/���H�.�y9�!O�����xhQǲ��t�ڻ��"�3	�B@e۬���Geڪ�Z�?{I�/(�PO���g~\0;;K��L������ ��d��	*�6�h{2�����dH�RY^6���;@v$�+`,��(a�t
+�Uw�"����[�!t�d�~{��r�f`����_[�5����چN�4ЁHC���=���U.��2݉��'��PQ(F��N��4'Yȱ�.Em��&#�R�j����<�}��$�ߗ%���妴ۏ�#�����Pz�Ms��9�� ���� XŸ�)Q��{�������c�W
��f-t���ٰ.���H��>[��LY�Һ�?��^�Iφz�gR9m�Yu4���7��D��0����-YnNP�|`��@���	Hz���)u��գc�T�t��|�R`I��uI�!w+A�O���������G�aI�p)`����E�
~�ь���IFs ����h�jw����0��[Zo`��]�20��7"c)l=��*t�Ø5T:��~?]��r��/�s�i�mu�G��JE�Q��0�����������\�p�OUժ.Uޱ?���I������#�*9 w�W�����%�k�ͪzP���%Rx
,�]7��u9�?���r�FU�>�ZM�h�������i�Z 1�7��
T2O�l^4���Q� �W��Xs���`�4��'�dɁ���2;mB2�x4أ���|��L3�F�1�_}�ojA�r��Xeғ�(Px��	�Z�m������?���ߩ��x.v�z ��qpd�'�rv�&����I"�L�4�t!����(�Xp�ͻ  I� ܨ��8ԊQz+��b]�X&���2��J���e��4sG��?�=������!j�M�OĮfUp��&g�jx���Go�@�b��W
)�$lT<&��;	$�i�{s�&�iN"�:��[����4�s�ӯ��w	C��7�h<�?U�V�Ω���b�Oh��՞Wl1�&A۝�f�촛Sh\[Yx�ai,�$���2Ծ3���A�@d1��E�;䠄�{!�#�T!���I=���2\4H�	0Pj�rPlݩwʓ'����fS:w��l�l��p��S���Gu_�ڹ!գ{�t�.��EO��T~Y�P0�HH�W��ǡ��`�g�lF�r�����qٯa1�k3.�cK�R�p���J���J�P�-�4vU���T���\7Gx�/�^�J�&��S7j
��$�?�'2����n���P	%��fnV�U�X�Q�*�{�ݧ�04\3���8Y ����u/e֌�Ng��_�T��aW>��
��ߵ=��j���r�tC�ө#��=�qD��B��|�.�SVWJ]�5,����U�cnY:��1���e�n��D�h��m��:��6U�n_�9z�s5�X��QJ��2k����9�r>L���c�,��a�ҖnG�d#��ֵ�)���cB�C7Rg2{U�@Ӣ��p�C	������"_Xsz��Bc�^Z�Emf��H�SV��b�a�K���-�Q Kȥg=�Mbl�_?�I�	8��v��D������}
���7 -̙��3����u�_���V��D�>y����+!�q��
�**T5<;��Y����]DW��� mM���La{�W7�%g����=�q$E�:ѱ
�B�~���r⊮�2�����>㇠[$�X(u(T�ż�mD����HPr��~��U}�w���m?�� �Y73��>x"�Prg�%�� ][��P���jmk=�NV���;�0��V��oGw�j����Ѐ��L*5��ʶD�!���7z�.C�X w|l�~�r\�v�2I��,�3OB	���4ޤ `��?�[|�EKm|ї�Vc��>���<�`՗� 61��l�q�L�L �-`�2�7��6@s`3�<n �̰�$#bQ��T�(c�癜�C0<���=�1��B6q�T1u�'$�:�'�/��Q���4uc�r� �7h���FBk|�kX��	0�O'�f�YƂ��F��yJ9{x�2�R��I2�^�=�7o�!s~�mW��^"�6Y�v�u��J��T!єk>|�k=�?��mji�hg��ꡚ��R� �*� r�q�F�N!��0|8$Ϳ)Q)�YL��'����J�F$W}�M�W��P���L���sܳ:I��x�濽E�qΕ9;��L�^u-��d��c*3y*�������r�z�,�E#'��V�&v�1Ҝn�Z�����k�{�{9S���e�]Re�7��3?��Ҹ�:����O _��/OO&���fx�Y��&l�9�it�NL�A��-�zX�\ۘ��If�<���Ox�"��4,aK��h���Z�J�M�N�,�/n�a��3#k<�W��ՊK��I��z���<�t5��!JT`�B�\#�_�d8��O#�� ���z��P%b�;��"z��4x��f�����)��>ٵ���f�X�Ɏ���>]M������kH�_C���l�o��P����n�y������{cP��A �C9�^�`���׵#��w�g}A"o�z�:Ԅ7K�����T�ף��i��P��*��Q> k���j\xG�����"Y�m=��U�4�5D����OG��.OW���ќS����nJPܞ?��^ˆ�"�O,��iM�~��9+��?)��8H�f��M'�-���5^��3ؕ�;]a�y%VI1�����ݡ|TȪl
�g	B��I(@ϵЅ':"*d�	w՟p��$�d��h�ud@�Fq~�S�?tD�q4���[�<���N��\��w?B��4�y��I`t#4�&{Oτʕ��%�]�nZjp�}��D6�,c���5�4k3���<HB��'�Þ�]}�%*�n,�)zZcX��;�p�������>U�Ё� i(O0��)p�6TT�	�a��e�(Ӻ��.��vvu���b�t�/HJ��r�%��N%Ă�ۊ%�Y�o�w������2i�.��Q�T�R*S�(���8Xގ��c_���TKO���znP�Q���:n�C�2 �M�!�dS�1��Q�{���p���דV�i��,`��5{���#-���QKnBmqn ���á	��BD�|�*l!#R��k�&���E�=h�Q�����R +�	��d\�o��F3G�|̶s�K�7%/�곝���@Fک�K�fH�ӂ&��sh wX�ų1;qةw8E��7T+L�Q.`�լb'����������n�)���ip�c����AGW$k)YX�l�%H[���^�Âdzm�EGݻ�υ:5YH7�e�1�C���Sl�Q��<ִ
8iX��z�i���eK7�R4�+mX3�L�7� �~]��Ԏ	�����p�S�ա�~r��Lk��<��\�$��!�X9��/O�sUR��=�YD�v(p�;�!m>&���&eC�x/sua7U���X�g���hwEk1�mlv��F�����?���� 	���^k���n¢�Q���ɹ@��P&4N\���(q�W�
�ڝ��M��zQ�FsjAW6NB*��&�}ϝ�S���%Q�c��%�-_�~Q�O��\��T�J��L�,�tv����}�~7k͓�җ-��j������/��<�h�1�5M�u y�:G&m�- �~��w�-��J�p��s��?J;6}��T|i��'$����"]	3i'��6�s��.D��U���M�5g� �{^�jč��F�4�~�ߦ��t�{���Ϟ��tM4S��W^Ur���s;|��}o�1������\s.����_���Y���Ju �!�xx�3/�"gg"�٬��s�x�7p��g|�~���Hx]Z�@ze����6'bw�-V���q�� ���/Y^�	IM⺃,:����&��/.	Pb�x� J?f@��C$sJ�0�Y�6J���8������Ae	Ѿ�1�J�Iͦ�� �I�[k���u)s4��+$�D�	#]��*�w��;4A((����9,�퀢v�����3�GHr�5`u�<֞��:��7�����r�=�0����$�d����������b��W��0�u!���@6�k�74�]�T�<A|e��Z�1f�N�Kya�F�b�h/&`�B`�n:`b�٣R�ţì���j>�B���5X�r�<�GF|]6B�s@~�(z��gY����	?�8g<�(Eғ�F�A3&~K	
Ŷ�'uF�s
��d��γ�nq�JlmO�v
�L�����D��]�a���w�W�?$���x��p��IPW���I�tu�4���X�F>�k7�)�}p[���*����d��Ң/P�{6�h��҈(V5�4 4&Hb����Iz��H��!�,s[M�����'6-��������������"�������}y��$������cba����R��yq8�:��G��w����7�!�!�:A%�0�������ox�NX�����_G��g��Ԇ��9n;J�B�͎�!9#��t�{~r�,���h��h��t2��v�RB�]���Z�V��U��)2�DvxHU�2#�(�K�e��v^�-�ZRB̅�� m��v�nj4@��%٢w�6D�F�^�0���F@�"]�U���)5��<1���{���/:4ӳ\���rt�^�E1��9+_H<�37�PZ����A"��E��D9r�����w�}�#PjS�.�R!TV�^y\����OW�U�.�,
>e殒�~��'�:}_�82�bN����aC���GۛGTA>671Q��D�����Wk�^�F-Em\�X&���@ٕ��T�Z�Nz-��]T.���X8m��UŐ���,��_Xy��u��V�Ѩ��/����*������L�R�/��߁I�۷�-�	��R��~� =��_
�)5��I]��R:#��@�Cf��W���p�7�<�|���%`>�TnDC]��7bY�*��6�>�0���n���~s�v��"�����8� �U�M���5�`�q��3��� s�3ݐH|��&۔R &D�j�B���|�]4JF��jB����Xs�1$�ܳ �=����!�:,:7��v�<XT8E����X.>��!r������i���9���/���ߦ�¦�^)^�+� ��U�0?	��@B[J�4�?��c�'����q�j�Oa(f��V���~m�q�b�i��O!gv�zo� ��Bݖtr�ؾ^����f�W�H/�>]:Ӓ9�t�[�B^0�<W��˵�Ո���c�w>�D7���3d]�P�6)F`��ΑȢ� x��2���<�
���
!i;��6��넃ƉL���98y����k�xnK.����F�C
��t�H=*�^��kW�l��{��H=�.�]AA���o��.=(�P�-}C�Zi!F��ǳ��5.GC����s��,��C������YP����E(�P��#?dg��l7���P�J~���L︓�qȱ��8�:�ڮ�>�dp�c_ꄶ+"kϚj+r���֔����Hڏ]0�5:�ʾ��ʏ�m��wG19~������ϕD��!�\n%�jX����M)|&_~��xMUrMI�Gʗ�le�!��g�[e�@�_�S���w[�W(�I���	�C�S���Ki�TT������Ǩ!���Z���+~�*����+���>ݥ���[B9/*�{КŢ��F"��27&��
{+�f����5~K�{!T��Pa�QĕA��2�h���m��ܠ/���PW�w�өS���-�����ݬ�ra8���$'o����X����A��2۸���>�,m���m%q��P���ۿ��R?��qn��*{ͨ�(���W���J��mH%�tƄc���Ct}^)g����̃ؖ�ڇ�>,d��=������a����m;?�Z���mN�+�[16V5�7o5�e��km��ߎ�L(��yJ�q`ylȴ�<d	�!���{=!H�+���x��޹�Z��^�/�N?$�)\D��SA�!��iB��������O#z��!���B ߙa�-��^�4�g��`� �ZqVj�+`�1��c$�g?��T��i�EU��o�"Ƚo<��;:?.�󠠮5��%���O^�8x�q�f�ߘ^>U�jE�_���槗�R�|�����m��P*'�p�j��z����F��-<5!��څ���ܽ��m)��!2���K0��h'f2"�S�\=+%ƺ턗��"5V�b����r�Z�z\���z�.���<�f�����oʜ,����ӿ�-珞��6K�( �h�t���lUE^�,*g֊dA���rc�������K��k�,��#�g���9�_l�!p�H0]��Vd�0��5�l�}Y�1��	S*-����w@�:�^�$IC�k'/�cJ4')ۘM7��8&�V�PFTw��o(`���2̮�=v�YQ=|Q�@�ȯD�K/	�ʏ��-�Vىۨ켸�����Hui塇4��e�� v����JQ7�qi0`���1pV��>�e7��L�U黍1Z ���5>a�����ț�B�W-��b�$V1��˚Dv ��:����h�;L����w ٨�&�z5��r��([RӿÖ~��Ij��ɇA�[�m�*�@�$K����)�h�'��s
�@�9� P�P�
d;E?Ѥ���������F�8?9}��͊���� �����2�[;n�`�+:��75��*��˧ C��B����Z��"���2`B���-�������_II�>ª?:<��IJ[����a�/	���QY�3�f�p>T��y^�ů�%���I^�8$��a�%���t�Uz�K���U5��Mv�R�sK@|Ub�Ң���5'��������3}�D{>sgy��vtF*XP��׈��*+�x�"U1���vb1�Β�����V0����,���3�%����)zh��i�Y�DՃ'��#��o�?�^��2�^"�Z�2	ǐaR[Ϡ�M!����7���*#X0��=\"<����y&�CVJ�*��x��g�ҷ����9�������K��2���@����`.���t�!\JyȜ�<0G�_��νlu��5�׌�K�5�4J�Bf�����p�{+����a����B�U��w>�&���k���+�â��ߊ���h�5��D�P<���O/6EM꫋��ЉOK�SCb��#��?�X�r7�B4��'ʦ1zߎY��7�{�8�t/S6CH^
�5 i�"��G�˅�&0j8�{!<�Z� h�+�э{� �Jp�绁��J�6fL
.l$�ܫ�f��G�`���y��(q�l�����f�0�v��IH2N��̒q7&Q�i�%5�����u��S�j*�����Jz�D	X��bmq/��ce0�j6��}l}��f��6<�����FM�|3[�,�]���G�c�vK��_7zb;�#����B7���~�WzDɱCp}�7\���<��}�F���E5@�8�iW�VX��_Pf����՟z	5H;F�"�X��C���5����fF�Ѕ�l{)JDƉ'V%sV+4��R؝s�f�8��J�=٥�YT�nb@@�k���X0?tD�\ʹ���Jq��Z(P�����9-��\���eI��������e�H�b���@!y�t�P\ϗF\��s��R���a�rw8�6yKhk��������rx�4��3
��{9�fC"�ϒ�����~ا45���my�1����s���+b�bFGm��_0��`;9���;1Gi�M��v��=[aL�JG�+�(��V��y��q�6CN��H�m�H�r{�v˹A�{�>j�yz�E��࿔��\<ԥ�ۋ5Z��8�?�!�F�-�C��r ���R��҃}��%"$��q��뫳�i��	�so�o�g�Y��0P�Y=�Ey-�z	"��}׈��%��KJ2N�L�9T�!��e�V���Vt��TOrTۇbAi8������S����M��C���P����9�醴��[L��"HG,2����W����\h�0gj�Ӎ}�E�5�w~�Y�)i�]�-�O ����~cפ�g��!R��b����,��,�����~M�뉠�0�a��d	�����!�}҃E@B����d��~��A1�x�=�w\��ǘEӋ�h�.@�y,�!�}x9�o/��w^�����p�T[���ȏ}���S٨"⡒a�Um3}{���8��4���6�h9�3�]y��И���tD�3�u%��q9�W�̙��Y��b9�e���X�c����1y���c/6�; ���5ޝXK��b�<�q�>�sG���%YG�_o%���A�Ցd�ot�~'�h'mZ����\l>��*A�yz2�nء��a��0J cH�	���k=+2�@Õm�t����%���Z��+ۚ�o��#�v /���o
�p��+o!���z��Ϯ����S�=oa/2�|�^�w��R��Z�����
H4DimDl!K����9����lVH~�d��#D�륔%�]P����p��c��½&<q��	�OZ=U[������E���:E�68fz��+�]c�e�L���_���D�u�
|晋�ߚ'�F��J�Ի�{��wWߘ����ao�/$a��6�nVps~'%��n"�)'�e���J��kC!�a�G�ʍ �?d�a*N�D��~F��z/�Q�z�:I+
:���#�AfE��mB���E�K�k���M��
H��X��/U��ȥ~;��N��Q�)��I�W����&�(;�ұ؆,�a�q=!��sԥ��� s/7��SA�S�	>�㨝ƨ�ȯ:\�&�=2]��!���kǯ4y=n�v!��xo���sٹ�0�(�@��uj�����6�FWk�r*N��1),�zI����^�R��x�ɓ�8M�rv��V:�w��0�]%>��xb��PR��}�L_�hd�<|�{��@��T�W���*�A] ����3Ý<�Z�h�G��۠"$���3Ӵ��GW8=m��(z��E��.u���N��دFZ�I�����Xq]�羸�����K+©�-�XO�a��y':���у:�`,��?v+�-�m��Ś�r%��`r�=��p)
�����f�6�?ܫ�"��8��\��3aW	��!/�)p���)Q��9�7�$��4�& E��J�UbPlX�h��`��l	J;X������X�͆���]ủ�����sc�"���P[�ݥܧ�1��|�$�﷉y����D�� ���O��?��C����}EqV��RraJ�~3���������V�:��׏���/��9AW�p������=R�.�W�ы��S�S"��CFD�b6̙oo,��!��N�����8��O.\�0��L�@ݪgd�Aq���g��R� o���Z	�#~���Y�*z��eێ��/'g5`�&]m�	����OT6�`$*W|$�;��o��5�2�!��j��D��L���ݠ˗x�@�nj���^�y����3S��Aoe�0Ys?���$v��h�v�	�<�Xp-���&5n��΂��Wn�]��ɽt�F dvb����p��D�yL�.\��4��4cj�LEx�e�ݟ`�%T��6�-�G�)��\�z/��zo���Z�aU%Һ/Z�u|[`A؏�cN=��^x�Z8#g�Md<d�8�H�I�/���j=\��rĩm<8Z�E�x	��7x���컞�@�x�s��DOQ1����K����4��:H:WcK�1Q���N���^yX#<��:-V�
�ڨ�X!��Q-U�w3U���ʅ�<g�D�8<���J���)�3M�6塥�Qw��$D-o<���=���-���B�[�A��d�{��L�Ok�olPk���r�
�Z����L�ET%�p��$��;�}�2��3NX���8VYyJ�!�ĺ&c�q��}ũ�?�	��,�ȏ�^$�+	�\[^ 5r+��=����ko�N:���hb0Mі̫����*\�#���<_ /�&Ը�	�������4"�Y������δ�k�;^�Ǯ5���@��dO��j�б��bfc�8���^��M�}��aU�I��(��X���"�zr���cP��6�.s��S���c�E$�f�j�����|9g�Uj�$��(�<QA��nF�_�7L���bf�;H����+9�f�2>�.2�1�8����-@
�5-�IxW.�Ԋ�v\�|�������f(����V����p�>y1��u�B�5�$�w��O�j�rN��AV�2���۞
�G/�6��a������OY������Y�kCdw:3k��	�!ڽ���Q}����֚"��l-Ax�z��dlB�	���Ĝ�Pq���R��۽jfD͙H�Z�x0�e��%�s:�c��c�T��ƍ���S��d�.�dD-zy^Lͮ��#+���Zi��:���9�f�� �>��P�j"�����y�L}wX���Ny�(����*Y��G�8%���|��R�	נ!����"�,g�>۶�v0	Db�����uɖ>'�x���]��m�ܦ@�p2v�|���]l� �x5����р�H��5�}*Y��s��2�������}�c�Z�K���NM78:��^T��in�9�_eiP���_��5�4�`�$���Wj0�N� �L>���pF�!�i�)C������-X	�풏�P�_�O��Z)(/�u]�X]�X}�JЄ�P����б�/�#B%�&@q�+�kU��ɝ��a��a��:|��&�_�El�%-�� ��Ju�{휥��;�W�VH��|ϩ��d�X9�LD��r�S��H`����uEfm>$K-�oH��z��R�׻��,��)ւ�!q��qc�]9�kX��P��C<���]4��0N�L���6bb�q�����C?}�p��I8p������Yj�c~�� 
Md�YNV�B��9���������tA��Y���	b;JPl�8����t���޾�0��/KԹ�k��0�9�k�>+�74f҆�\�`v�$��\��Y��O_��H��F�r��{8�DK���_������*v�T��Zx!.V�I�B���Ķ������z�R������"{�P��H�?!O���k� �ܒ��gϯ%��}�d��a	����S�N��FkN W��×S\Di�S�Bc>d�m/�*�Gc���"vZkXr+�)-S�k1��8m�����W�r=���<q��ڃ�܏�9��`�Ч��$A/��ذ��D�2e��n��ٕ�t|�ﶶZ䥬g?Ő�b�6�HN��Ρ��(j�Q�#�&�	�A*���<]+��Bz_��/׸�݀�i0����ه�J�:���f�����x��,�S
3�C5�y�*���;�F��M����U�a�,j�d���a�"���n]c�~�#�pX%#.o������������.�4�[���6�0�@n�yL�-�O=�s}�T�PR"�"㒲g���H����$�1���17�o��x�N�vF��e�ck1�J��ҽA������_�m37Z�O;~���~"$	\���S��="��Ut8�L��'���J@����G��JҌ0���?�5��EHn�l?#>�����¬7��g:� ��0x��Ю/Û��e�d7f�.I2[?�i�`�A���	�s�À���e�u�OQ�(��e�����x2#=�Y�t~\K������S~����!�#�7L����X!�0�o���&�I��d�	�*���6���8Ub@fO�wlu��=�Tsݮ�Vg��]�"�7#�s7�R5���6%ԒyT8�Ght���g�l�L-��+�ɘ�@*El]��D���G�=�`^oq��ť�2�����z�a�UR����"�GD�C@y�&4�V��GR4��h�	y��T	.FZ"��\��l&4�n@��������e1��5B��v}�j�7��A��!/y���'�F�Ғ�r-�RZ� ��w@Ͻ�-��"����%g����@"H���Puݠ�!���̗��Δ_��f��9��v����Z�Tf��u�ϗOpd��.y���m�f`k]���*D�S�������
��M��rL��묪����^���z+�m�ǀ��6��+��\@�S����`�˨ݻJ;�W�S<�R�󛵝�r����̥�C��
��r�"��⡅�_=V�zN������ޕ~;�/|DL�M�}й#}E��	屻����q[�O"#����3��L�!��h��a~US��#X��נr7�<���˼�lf?}LK�ԓ)���( �wE�B̽&�>î��[ ��-�cĐ�S�:^UE�*&�F��F>�r�\�~�;�ɔ�������<H��Tm��a���Ok���^o:��se������G������Y27c��k��P�&�]�4���.����a{�F$��=����~�C�z5.�r�`�AJ��8p�δ���M�#���˝��9T���7�33s��a���w����Z_!�l�a;偛57Y�~�lG��1������-�����\�F��#�G�u�Cqg� SE�����2n,/���V�ɶ�����E)�]FA���)ļհI��
��$��u'�)�S�Q��������W�H��w���W��g\�i-�	ȝ6�|�6��pn.����Jns�PX�Z�YG�Q\b)ww\<����R~��v�������x5 ���n��N�� ��-śM!���Z�p�6�CDp�`�K�S.
 2H$rU���́H��j^AR����0;�V�UI m��lZ�?�f%a҂�L��x:� ��K��4��x�S�3#�@,T捖�y�X���4˘EZٻom6؂o���BF{�!�Xm��-d^�C�V�¯�Ī�tWh��4�����^��q��lUg�[�E� +�Zi�a����8_o�w���7�z�� y���_+v�j�����]%�tx�7v�z�|lS��|�v����q���*�+�va�h�f����G&Q�ȸ񆅑ઔr<J�M]��(z�~����X-H��@�o$W��kxo�0^B�Z�e�SӠ�#�G.9���ǎ��	9Q�w�����[�Ơ��&��`B�3�9G>������M����h4G�/׿f��(�DB+ɐ��~�24�Ϡu�
T�^4fpE$p���hP�x�T�6�+��,�/պ�b�����_l��(���aM���!S:��S���ُ��d��$W���4E�q�� ל��=e�E8�d�Ru���K T����~� n�9[�k!���1�B��Y�1���͗��ƕW��h�`�(�J+b�����1��3>��e�O$y2��N5!�Y�G�6#H�&�0C+�]g�N�$�"w._�����R�Y��@�;�j�,z���~ppY��/0u Xإ7p��L~�6sĽ��+2�qx��u��������&(�
2�)\��D9�p}�X����jSS�o�^�$;X���n*$���7#z�n��f^�� �_A�/R4����"�U���;R7rNhі����ظR_/'�'�XÕ߹��Ѫ"W��g����>��sͮ�)�ޗNQ,i���dbo�����M�d���X��ko]�F��gQu_R���P�W�3��Q�s��R��&9���R��cP����t\�o˟w�8-།��.���[e]�4�"��'ʨ�p�$S���e�F���w������BpVS�wpaQM�������F��8�)��g�p!"�筭*#���ı7��6�.�H�'ưY� N�C�/:������ 2%&���ijᘥ���Py�d�d�iG�_�+����˷�r~�-s��A����b��6���{�~����<�ha�Ӛ�n���R���ވ�N��B	��e kp~@�Sd�S�M��j�2J�,qf#�q���� �&�� 7�&�B�N~�ײ�$���>}�C����j�}YЃ|E�scKی#�!5GZON#'���P�q��I�OJ`��A�"-���0It7�30�Άy$��Y6	�\�L��d�O֔�9���n>9��'	�SX��Y
�D�⍸�h��̄|�����m|f�:��>�����%�� yJ�
��~�K}7l>��;1?GLUt��.��G5�6�OH�2���̭�B�hK�ë�O�<��7��U=9�ӗ�޷X85I�������$�D���(Яc�#X��S���kA� g�ͥ=CrW�Z:T�Z��M&��5��M�8����%2C�i���"+?��v+ԃ���O�o��9�?�^�;�I{��\�oݡ�w)�41O�B�<��
��ɕh�J���q�M�������x��Dۚ�h�� ���K��8,෱��]�����r��s˲�P���	�������D�Q�L�	;�8�:cVk[j=F8g-��䘽j�X����vf��5;ۦ�P�Q�D�V����p��X�-��Nu��<
ەW;/�WB��*�v�&��ͳO�� k,+�����7����m5��V���(\��h\T?��K�8ͮ�(`K��������P>xr6��_�thy473�x�a+�^��H�O@�;"��`��E�s����H�
�SF�{���!@�v��~��_�,�
2(l�Fw�K`w+��z,�߹��G��GZ�("���p������ihP��O�ZȮ�I�������|�L���n!о�5{� �oGx����n31\����~���{Q˪ �n�����_�P�ވ��՜A�+���!4ۅ1��S��GP9&�F�_�EZƎ�R�r���>ob��FQ����8={�c}�ԃի���m^>�hg,�4�Y�^pR�a��j�mϜm\l���%�3��Y�8������X�\���'�F2D�� ��D��g+�9�R1�P�p�#�A���}c��E��3����==פf����7R=��kޓ|ct?HV�3k��}ʆ�������E"x
N����4�Z[~he,�����P*-���`�$���
	�t��g�rh�k���]���Z��̢��ޣ}Mޫ�*�E��LX�[ȔY?��:\���B{�N4��[���)�P���t� �8\2��-�핞�_��� �))�F��7�`p����ಳcRqr ?�oQvt5��4����C��c'z���jy�U��P�$K �u���4e�@Ĕ,��p�P�EƦ���=�n1LEH�a��=���+�`I��bW�n�*�e��G���I �6�O'�9B��?㰠{�n�Z-�M���[��k���).�;2�\����Ȑ0�22�%���kBU�2�b�8�r���Q�IͰk�<:��Ng(���x���?�΂g��v3�R���ev̮=����A�e㉩O�jO����*PyD)�]D<�Rr�qT�Cv</����Q��Dk����B�X%<,M���R����?Sr&��	M0XLk*���m�����-
�@}��<�+��cf+��Kp�[�L��_1{��+�T)_����޼X�LY���-Um3�0���S��g�luqF �X����O�d�=����Lbc�Kkr��OLH���|�5�Z΁����=���$R����:�Y������N�Ű>,pF
z��JR���E��^l�"f�]C�rcAL���k���[��Z��D�Y*�DZB���@�6r�`z+/����*� #m��W�V������Q�eF��U�&ˑ����C�R3c�m��O���-�s��ܶ.�9�hI0AV�70V���S����M����X�+�h��C�m.���Q��R�+#;�Q6ï�^B�y�$��$f��?c�x��������V�#�۵O
f�}�iR'��Ǘ�n�`N�|5Gm�fX��8���X�|}�q'�����˸� س���]�C
Z��>�9�ɚ!�aO!�ue�n���U׊Hv�Efa�3�{#.���Sb�qǀ`I
!�:���i�h�#����ZNd�����Rn+�
�ڌ���(�+����y
�%">Fy��t�7H����*�ίT5ʋ�2����"}�T�0�/�i=V���q9���ku�Ot+c���w��q��S3vg������@}�6s��`�W$	\�,���K!OX����6��݋��A+����(B��D8�L�*&=������5`� K{����@�A�A�.Վ���Q���`v�Tπ�݆`��%6��.�
a6@�N���"j��K�?���åu��|I�^6���9L������{������k���|�5��J)1|�p��������6���ό}��x5�@م2� �h�{�r�A>U�D(�L�𮮀�!B����mKfߓ���� @/�k�Y�����������U��_�P
�-�eB��'j��e]k>���\ 31Ҩ Ĵ�f"���Kc3���~KBE3�6�~r�^0�QҜ��c����~{�e���R0����`|���wv�VV���i�w�1[�ګ��å�q�7������e�^W^�p���uq�������f�/Q>=3^�;�̖�E�N�t����0g��8쫾��	1��nD�O=�W�� ��MZBOw�� �'����Rh;�\~T�N���m��&-��i$O+�\��MZ⫱���D�Wa�"�3��zFU����������e�=35�6��n��Xo�Xa�>��ٯ~SjU?����֛�����b#IϾ���6�[��<��`f"��]୆$��H�/ g���{ Sc��vժ�ed�ٴ�j�q�[��.86x��?c��Mŧ�A�9P�m�GO��>�;�ǌ��7�V��/����zg��������_�}P�[Y�g�������� S�rX��@:���X�$����铊��͑r�̳q3y����HCLa=��$'2�hi����g��8�*�E�oZ���6��5��8
7yp,H�7�������>�A�&<z|n���m'Re�S12��@@͞�p�d`�F���%V���%�T�U�!3������DmoV��c��&h��;��S��د��)z��T�-��p)�)(f�����7$���9$��"��@o�	�p�{�DZYa��x�i�k-�]|�%��IJ)i�p�2!J@��zkI*���_�*���Ȯ.2[����qY�1�c�`������e]M\Ї�l��Dю���:��vv��'q{����c�>��t��I$�����	��c�{�����3?Zn��,�N�(UW���W��ү��՜o�ܩg�����#��@�F\$ED��,V���2����i��f��6�з"����P�?�B���Yl3P/9Z��{���S���>������!Z�Z��������;�y�v��s�3�"H��+VL�G�tM=�نHM	�-LP:���oQ.�tKۯ����5	��v 6LJ��!_�qHd?��� !�j�A��F��o\���h�Pg}WL��?0������y���G_:\� � 'n�~��њ[R��hǈ�|�.��2���E)�s�?�\���*ƿ����*�~?�,��A�Ǒ���!��AC�_��5W�v��{KK�1�1���!����3����Ϸ����c�Px=�����7��rk�[���5���#2��~�c���V�c5A���Z�=	�q���`�3��q�8R_[��b�۴��6p��>�*Rq;��/�6�jI�i��)&r�ru�]$t�m�o���u6���{<mÉ�Y���>��S�
@�}�1)�#A�|%"�ɢ0�ߚ�2D���B��y@R�Q��/L�P]�	#�S�s(�=��tL��H�8ٙ1d��rJ������zO�
U'A��q�'n� ~PŨ��;�{�
&J�ŗh�ᬐ��K�J��c���f>��=�B�ݺ+o�H|�2
ً����-�N��*������6_�L��i+�6=�s�g<As�n��B��qCM?x��兑����Al(�*0�T,�(yu=��ζ�b���׌A�� �`c�ߤhm���;�6�����%����qS�4�?H�_�ɥ\�겘��;����Ss�Y4�S�(J&��Y`���d����-]Ҳ��5qDadY�p�1��Y�����5��T�A��'I	́2'�J��a�(n�ݰnv����H4�@�5�&i���&��_e�낑��Ǜ��F������6gI�+�ۋ���'�;$��/~eHL lc(nggj��t����F�hh]��9]���"�{]H�^w���!�C�7��W�׽�3���t�]��>:6㗶����FD�4�kE5n�ʳp��i���e�]�r�����e-�=�ŘQ���SB���L^%��k�7T+ߜ�+����]؄b���8�i��L_$�l�0	��ҳ/b�����Ȏ���֔5� sv5~�D󠳽b3�����;j�ܵ�- �B/OT2�>����/���\*B\-M�L1,9e�FX)�cC�Ǣ1e�o��'�-wǖo��`�f��6u+�V��Hm�)��Il��X�ev�8Y5q� r6��D�z4nD��UZL�5��[	;
��tO���:��bx��C���\�﨤S�ӹ�|?Fs�L\�'��F�)��P���R��I��ꣃ�����6R�������W����
[A6�CUH��;�f��E��7¢�^&MyJ�N��ai�ۢa߰#H�o%��&���sfo��A��rfv5>s΃,����V=�w��nErL�2GۗU�&��\�-4'=1�Xr�އ��h�3*Ysê{��& Hw��0�7���x3�4�p����*8��u+������h����W��Jyp��)E��s8�EV�Y�\v
}u�	�N���wBS+��HH�� �/��U�/
�P4���H���ƣj�'����{,w��}�zC������; �*��|��Ý0 �񧎖�:Zv���'��B��5tw�D�(��Õ�k���L���ٯ�O�L�3B�}|w�B�;݅�]0��9k���[P)�<�I��h:e��	�T��uUS0Q�I��a�x�||S1�*��a�'�(:��Ÿ}�2RQ�C�
�zq��5Q�[���||�iՍǴ�7)�0"FI;�����^�1��H��$��2���]_6[9z+�F=@Yj MQ��~�����cn�o�>s�_��0[O��n�B��[{J2hym��Ѻ,n;�-I�L�����D��TMߡ��Ԇй��ow���F/SC���C/��I����5���־�Ć�N�	�(׋�lZw}����B��ިl��d��*��L�.���q�
%W<{��b���}h�T'�,x2���qs����D��|p�ӽ�߭FHc�<ˋ����m.
{-fVRfC\��[�Cv�>93��9�	��?RQ?OPT�%z_+)![�3�$j�*��w��ސ��dB�m��B �����]��]�x��Nh$���l���P����$�+v�3@���7	f�U��-�y��T}y���<���S��8�L�逝��}P'�R9��͈/��VE����`����dg�ǔ/v[�=am�z�G(1�&��s�)w�/�<r�F�bntX���K�� �ˊ~6�������"�����C����UP��V�{Y�q��E�	V�xzhN���-6�6�␽�X�8T�U!���cN���o唉��O �3	��(�l����Ӕz�dεyC���.�` 9H_�����5��D4&�r��lɵ��٣��H`�bR�%��;9��r�(gم;��g�Y{�F�_I=OH�vq��������rR=��4�]�ʚ���̿����,sۙ���b\=�}�-��j��+hy�UpL� [�(%�ёCA�;J'T߱��$Y�`�σ�(fT�6pA���?������&�Kp8vk A��� �ʓx�X�<Tm���`U" ,�x
���������:b.}@�C�rFe�k���[��I�f&��5�L��-i��85C��A�o��9�y��)���5a:�@�h����E���Q		ZzQ�[�����9co7��/�\r�4Y�#7�>��\�An��yۻ�g�O8e)����Po;IuAv#��=�'D@��q�S��7#	��N=ּ��Û���h�2N+�u�w��L��;Lᵿ�i4nǣ�O%ףހC�nӘ���DD8�!B*���K1)��/k
�Դkt?"�I��g.��I��P��	Z@��'+G'���F�ђ����G��30Q,���3��7t���#��J�RW�:w� >�z�,r��EF��k�)~�BiN/�M�P�{]�sT%������F<��Q�)��.��b�-
��C0�����	�KAAQO��j<PB[�G�v�, y���q�H�Ӿ��q?,��*�����w=�n���
 V3�xwj//�)�I���{rK��\SV��J�Vʤ�9��0�|jt�ɣ�`��!$/[��%"�x	��G��M��2��T06���կ�gh����6O.��q�Oʙr���9�(��j�+_�q��z�Ǯ��X���̫�(X!�b�'*Uf��#�qh'	a�l@XV'��0��M�ɛ���ȇXJ+v�}T�x:�D�V��h��̳���v�,��$R�K���a�Jqy#�9H���h��.48B���_p6��Wj�$�mG�ڴl4(n�aon#�PHOqK�%Pj5��#���Ͳkl��F�nKi	��I�#�J�[{�z��3��y�mLҐ'�ëд)v���xڷRLP?����$���?8Yj��w��љ��X~�� ;�:��V�L\�$D����qc�v�uyY�7�\È��`�� {KG��N]�<3���]��DH��=�Z+��c��56��^"�F����k���{7A�gV"w:��p�3�s��|S�|'�>��&+O3ى}��'Cxj'�?(gl��������my�� ��@�bG�TQ���g���<Sn=LoQ�q�'�NQ�M5[-�$��%�#t��]t���t/C��)�L=�w3a�1?�!�ܵaL���G&����A}D�d�� �ߎ��\��Q�,�uP����6rHJ_�����+��R �q/S	(�c����c��	E{à(��J)�����yh.��S�!��/��Mg����*y���g�M�vh	+7[ ��Ƅ#���o�̛��ז�UO�W:�Ȧ̚�!t��cm���ʤK,v������C ّ�Z���d/�F'.􍸹�@�D,�J+	=����D�{���Li��U���`^���R�1	��`��w��AaTdx���Ե[s�A1�W����A��w�]���k ���.�vq�����5��%�Ue�2����!vT$�Z����U�H����es�,z�,m:3��P��4u0��l�����n	���t�DWjN��Hf��%�>���э�%x�I����*Â��(�3��p���6D~W)_�y��=���Zr������s��쵕0ϼ�<]��i�d��C��ah_��#�S?o)�[��������,�*����̄>\h=U�r{yQ~��]�s|'�7����A.N��|��gK��C�`�j�4� ����dfn���6/�1��J{���xޥA��b��x�߄���3�Gq����&:(/Z�-�����M�:P/��N����2�E��L�V{�6o��hf���0knb'����W�-���>�
|��H��3:�3(C����b"�D�����υ�����]�!�'Qp��ʡQME���k�Q�Y8{J�ʟ��uK ���z��06[���I��� �	6&���J���ں��U4l�S�N�ǖ���w���6C�d�l�0B2�@?�L�$����W�v@���y�Q��-�ty�ГBQ��9���V���:v���CM���}So`��bS�g��dv���W�a��P�àt�Yx��ȅJ`}��$Ҋs��7����sMl�Ɋ�<�c=�<�afl��sd���>�v`��5\o�`�MGl~;��n��0��Ɠ�}"t-���=�+3\�&޲��=�&59j�v\��z��<��#i��9��k"���:�5Ѓ�)Rq��%�k��d�5Y(�>���X����:.�%2o���S��`��"i�D��c#@j,�`���^��~Ǫއk��D���"r��GP���>�N�W�b
�n��� V:�FK��%�8���,�Lݣ�I2�Z!	}�?�5J���g��ՕiԤ���Q�F:��F�-~X�	�5���,EU��P�)��!��b�(��QM��Z�\�;�6W�26==�8Z�7�v�q%����<�ՕzePONYE5:���7�8&�r�{�Г/��H��h>3�ĲX�U�S�2g�X�a�Tqv�'�����v�|�n�%c�Iy��e7����Qz3t�JH��B����ѵ�f֟��-�0�PB�s0��X:�����CEx�K���#�6�wA����y��I˔9��I����ߢ��n�C�J�����5�<���vyc�"~~�<���/��`~&�7<:��Xx�DZN;�^���?I�
D��9�Ci�j�����ޡ���z������z3׌(�/��h�~f�?��R��վʗ�>w�$�����k�>-g�J�L�����t���A<S�Z� v�l�c, t���:�3����I���3�'L�R̒-�a=��G�����A�|���f�ܯ�tj��)�~� ����H����q��V�J�+��Ҭȱc�M�y#4y'��;��R%�y%�[��Cǵ�2jn�j��-���#�Х�A�������%$"?L�I�hҧƱX�{�ݯcXc@��] 1�˓d��Dy� �*���x!��t��L�Õ+�}��?�߼����#��M���V�u���õFr�N���*�/�RST�J��6+۝[�=�]M!�L���@6{=
��A���H{��BD�i���|�/�[�B��)��R߬�U�-v$�*Wm��C3�-��z�X�A�� Q�[��U�F�m��RFHƢ���{/�T�����N�j���o�EiDڎ�%��		�r�B�h�H��R�(�9E"O�]�N�c��I�`nՍ{P2���b��B�ǹ�tћ����,c��P�'3Xŋ��,E�l���&[eed��5 ������*}��D�D;a��Q����e�ulЌsQa2E4�5}@�k��δDE-���c��WP�Y\F�6Be��h��wY[Ȑ~px���s�:{9ǅ}��Ai����ӷ��P�i�Li�t1ؠSH�tFԮssV�y逜Y7�.Έ.�D��;Ĝ��d��0���B�Y|O�'~�"���k`�`6�$����
`���d����3A]�6]�&ׁ�@��U�U5�B�I*��B��0�w�i���ٰm ��y��~ߐs`�x���� �~�-��nT�`^<c|,�$n&��Q5:���o~<N>Z/�R��t���'dZJ����kY���g�<���g��
)H	i-���l�.�]?~B}��w�X��lA�v�}��UV���-�؟���sk�"IǺc���J��z��:���<�>�fq��&���v$�XC��Q�2��41Y��y�H�5m�NȇS���NX@�4R�F�!��d�2���`}t�G�H�WΌ�=O] ��ғ�7HV��i�M�.J��_��c�m�
y�	���g�GE��x��u�XqB�v��J��ʏ��qU`���T��F� �g#+�+�EdP�E�Y#L�b�����R"qg��6���@�Y�|�g�V�� ��kDA� Ft�]��+��)ya���� ��N���ǊG�$��a6"|�x,��I�
����zW"���b�$G��O�#+F�8�l�pZ��L��xa-`�U��!�8���ka��Cc\@�na�-������g^�h�;ո��,���Tm8R��+d_9a�'d�� 'h]Ukg��5�YG|@�'�(���ҦO��'G�?q Ґ[�Ƿ ΍�����έ�~]n�UP��q���Y���9�	cԐ[��8�h����6�� O��
����)���2������}�yO�I����J�@{�r@�D}��n�s����@�66�L`�L'�[X�BP�.�0H�QW��l� �����u𫋨��mE��O�zbݯM��Ч1��+f̱!q��zTl(�J�k��r�@����D<YK�@�nC_N�}���-C���8���Ӌ틘R����ΐ�+��}%��M���/܊z��9KT���_f�G�d]�a�@g�{�z�3�r�!f�JP�5�����w m5RњL�,boOw����B�.����(v78�V$�����p>����1��N�� t��;4���r/��6�;��Q���!���6�و�\��R+]rF�c��	.�q^�eˢFH����9��L���M���*;��r�M�~	r�ě>rER�MgQ�Q��3�a���ll�X�Q�&�kC9�+�Y	�Y��=ĉ�nD�ee#W8��%{�X;=�~G��Z����NrQ�-�cG�=M�[;���ɘ�;���%w>��h�����6��H?� ��Y�p�
�}��a���wYR��g��Jy���3f��N�mّ~3�@��g �\�FZ����:�N�jfE��#��1R�Jxtk(!���KŞ��F�Ќ�lC�Z��X�wu���WH�{�e=�.�y0K�}�\Q��:��
���&Q%��
�p�H=gDZ�&�6�Z!3G��F0$�.p�E.Y=��_a�g)���a�M'�9r�N��ne�d)]�;#3��UG#�7�4�;FT-m�7�")@W� %+d�j���M�o��91|��2�G��/��|6H��:�+j��_(�Dϸ��'�!Muj	�g}̚LJ��C3|�y�Ҥ}�x�x8�>l��~�W,h�[g1�!r}��� �<(���`�is�倏f�xG#��_ �yQ���|x�D�xwePm�0��z.�l\)��	0���Op�~�cA�7�2&�Z܇�q\3�L���SA�"���Y��J�� �7��XC�?P+9	AȨ�^T/��pg-[��ȩ	�t�N�j�s�G\�� <����e�@�����g}?�-����<��l���v�?-�S�����Rq'��0_��� ֬~�s�.� ����;�$�!!g�vfQ���5�t3��ƒ���b�u�����&O�_�0ғ��ީF��������6k?u#	2��4��<a���;�5�t��Bi�3ڷ'��Twl7����d�XT,s&�z��g����1�Ei���% Go���k�9q,�o�~h�pkF������jը��K�K�=2�D�J���f��㥁.nwtk1�
��s��,�8&�a0`=����WE��w�2SpB��Ӷ7�57�2p�J�\��qs<ABm�	�,���Q�0j��Z����u��aF^VW��9v�.��ӯ�<�Ad�3�y>�s�����r^|�,��!��xk$$䝌+��O�(J�E�p�ԗ�c0��` G����a�؊'{���^��@�0���խ���X���)|3nl�B���$��]��o�3ZM�Xz��B�e�5��ʳ ѯ9��0&O�݋���B�:ǵ��Z�Fр�/[�1	����B�D߂��A�t^�jQ�3d�����#�el�iij�����f[2�5�������~b}$oiI�l��e6��P,Ol����dޡlg'��m�m�VކO�V`n�EhC����d�	,�s���@d�\���%��3��Db\Y|����/W��v[s�o+���t�����8�݈Ϛ�I��xƾ���c�����iS�������y/��߸>E��j�U��lv��4�˫fѾ�Pp��`赣���Ac��֤z��::ɐ7Ԏ��(����\U�S�AR�(����-�X*�)׉����U�LS=;9}�4�����6���V^����і���Ew�]]:uR���"�3�L��K�� g��,�>  (�R�J���a/?ܔ�u��x��#R��1�T��3�����i��ע3�Hn���&�!�M(:\�E���X^�:�4hu����F�S%,�jv� �A���`�?�x��}Nl=E�̞���B��H���Q!g���8N���_$鬅nK�&ป�4�k�X��I��xP���cr)r�i��C�����sӁ�]���.�h4�0Ʉ�7�'聍�T[t7*�t?�<�w���W�F�i������	�Yh��o[������[�����
�_�}����j"lE"4������1��wD�����4�Y2n���:.�c�[����)e����C��6��#]�;���m*�V��ee�ySe�G�f3;��T�j�"�j!�v`�G'�SF4-T�	 r<�9���&!$�t�}*ne\S"�y^�m=#b�/�Հ���$�r��(��+Ss�U=�-/�n'.������g����hKm��i����:��	j��0��Ry*Фp;�U	(���w������E�q�qa�M�����޺G9����[fv��蹎���N�w�f#�Ƭ�g�,�3�7�n{_����4���m����>LxQ9��ݳ�ddK췓P�e��p�XV��	3Z��x�������a���������*���hN|�c%\n�C&��fsSv�Ƞ�:F�9�����F���������QZ�~h�P����,��z�F8��,XYJ�ܖ�C��Se�X��[���KÅ���0�;�cGl���Ӂ��[�:���E���*0��sD�ǆ��1�����7�4�4��*��>�30��b���[7���T�4ȕ�j��=Yt>��'Zd�џ��t^�T�F[�;]�72W.|qJP+��r@l������N����r- h���T�uo�Q;Y�uc�׼�D��q�:���+Sm6J�r!j�m��)��֗�ϩ�1=��>:�ʳ;]�q
�3fr��^\7Պ���O�m��-B�7�4"���J��zUr�D*ʹ)-i <z�����6����;x+H#�2�l>:�+T�����>��1��nO0o��)qQ�`K�����q0���i�<o�rP�"��T~������'�q��s�P�2����"�_=�������t���P(�sls�:���)�!H˚�SkܛZ�؞} ��NP��J����m�Z���_/�n�������,7��R���ם\!Y�g�z�#w��5�������EU`�5�P��1��tOjb�̄�dd*�5���L�]nE��`'Nǲv&T<�x3d�|;IǺ��YMC�"�Y�����^��t������O�ĳ������n�k�b^��n/�:7)4�Dy*;z�bG�Q\C"j�?�����'(-��M������y&��_�^��?י˧�T���yX	ľEL@�����#n�M�M�q��}�&)�Dgl�c�����hU<���c�xS=�"oj�taϝ��^�ł�S��J7b�H:����bb�m�GbFD�n�k�=��3�y�)���wOJ�hU�$A��#�j���0�H�iY-�w����p}z��ʅ�\1]x�EfAy��cтg��c黢�ʀ�p���_	������G�# ^SL��t�x��!�-,�;�F�b���n����q�CY�-f�)���'���p�w7A�@��D5Su���p9��ڈЅ}<���J�X�����<8B4�\�wfY �)����p��z�;�Ĩ�<��+	j�5;7�K�h�i4��3郜��B�8x��>�*81�	R�r�̾�\Å����T���J�>MPƲz�1} N��iQ��^ޭ��\����8����3{Vv�q���ð'�d���6`��T=��31�_N����;�dyqX=�;�]��*�c� @��҅�4��f~�^��b�3�c�TB����R��ף?o�L�h�6��M�$yo++���D�⼟�h�����u�h?q�(¶�Xs �I#��|�[�Vư��%�~�:qvX[֩��T���j!5?�@���rp�n�Ƿ o�-5N�����l�A?�pZE��<�.zkI�@�%��\7^�>ck�w��F�Y��p�vA�}�L�G�3��tW�"��)Лr�GuFo���L�PUFO��n�A�@,�ڧ�B�W�so�0��];πXR��9�@��q��˘�˶d�ǔ_��x���џ�����2��������1�}&���heOɅH]KV�d��"�ի횰G��+k�#���zĄ��ы���Y��t�H�v��ޠ�v��V�h�]hԼ"
w%�*�|M��#g.�7a�$��w�[F�;���8�8li�]0�N��)��������W���XT�%��n�&�`卧r�a�gg����J����A��Pj��Ż�\��.�)��������h�IΨ��+����RM��g���8h�7����������̱Hf��cDg]�'U9n���:P�Y`B-ZQ��Y;G�%��eۮb_1u�"L����:���q
��>;�Ѹo������j�eu�R���'ޮ��6+Yc]qW�dC<K�|*wvʮ�G�L4,J�������M���X��Лg�_���OaLẜѥ`-�Թ�ĳ����Қ|�7�Q0�
���h]�n�K-�̣i`zc[@mT�Q��0��!P�މ�Z�~�Iެ�"��Ź�ص���ҩ߄����gͺ����_�l�
W�ن�Dg0��}���,���y��[�2p����g;����{a��P�y3\��-���gڵ������ڳ-؜s�=��X�6�w���c��A�*��� ����@&�
<2%]]���;��8��/�0.wY����"�n5�u��'���|=�:���a��e�Eܗ�xO�y�e"��8�8���5{b��TJ�#�G�����2f��mq�*���/ b�s�l�:�הσS�&8��.�E9�z�tX͜��`.$D%>����qh_�vpx�����������b\��Zb�9�m���Jm��t���l���� �Tk�B�D���9���j�}�]xF��)?q=ʵ1�J <�_aCf�Cx�qշ����N˃8��hr7�2�[�n$�'dL�ҟJj�򦙄�/J���,�4B���1CWu�A�u��$����L�O��`汧u�g��Uu�qב��]!��d`���n*"cG�d&�еD�Yl<��> #R����[2�G�D�`w�69�������8&z=�	�*���y@	.r/��8ֳ�c_Vx���T:�3:���&l�HY5u�*�W��^ɵA�jں��y�OET� ����ܻ�:���������bc�,N��h�RhT�!H�S�O��2��
��8:G�>åc��0���CD��d��.��:^Q:���H$�8���E�"�o�2�*wM�;9�s���<[{F��᡽���蘃��H��KȖ���4Tu�q�,}�`���J�xk6����Drr:��Q�$��E�/�0�g�~�A�x�8�}?����.��5ڜf���Ӷ��e ��Oc��ޱ��s��{a��o�V���ɱA�}��Z�7�j��=o��~bw2"�`t�O�t�d��vQ>�i�?H��
�z�w��ʏ�y�P��o��F1f/�YgnC�_�F�ۛ�ZW��A�C����D[��i��C�u�Z�i+�R�3�<�$Ť'ɼj�bhV4�m�i�}��00oT��i DV����&t5�'jܖO�Ķ�Q\ө�5�X3P��B��}��̾�u�֖g���۔AG­UyQPxN]�X6�9~`&�%[��8� Q��7�}������w���wC|��lJlxʧ�:�;���W��7��t_���H1�!9��yȔ�FsJ�I+&�Wp���w
�xA�9�º^����χʊB
�8��yƊ���k!�u�I����F�R<��=�m�<O�$O�˟��_T���T�:8d�F����͗B��Y��H[U+���9�9���p��������]1r��hlQ1Q/ױ�GǶ>�:���W?]���EI~�b"��8L�q�9��a��X0lW�oͦpf[JE4�Շ}(�91��Mژ���?&-	������~J�����\Tc[�6�B�<܇�D�B�9Vh�[����x�׳�/�g������~��@
�-��z�uUgY�ۭ��#�)_����E���
 щ��HI�5G$�*bpΦ$'��5Qg}HS��_E��CHŏ�)b_=L=��]ag�c�� � ��ۯ���{`+�Y�+%|��W��BGX�I����[_�uP�ڳ�&O�Z�f~ ۈ}V�T�.Z`:ZD�qE/���Qr�h�i�/�C"pټ ����_�v�
ŏ�F"ڒ�������k
�,�^S�����0�j��f��D�M�wE�֑�/(���T�x;хox��w�� R!`�}X����T�Da��?Q,�4���ڞ���]�%�������Ri�Az� ��{�����,=ķ��Y�PL2/�_&}��>����u��p��MKH���V�3�g7�Dl���У�b������a��{�4<t[�YuU6�=�Q��%`������{ap����"L��!l�$���(��.x���^���Ylp.E�M(Zfv> p��Y��ܿ9���T�s�a�[u���*�ͱ%�;:/if�5 �)bCy��/��P[�=��D'f�g\p����B�v��|V��{�o����{Řr�b���c�'%[�eb!����^�~�M^�EʩXW�WH���p������Z�n=�n=mv�X�R��D�@e;XA���͖5h������Ŷ����313�3�6�!�Ʉ0����*\z?$��|�{�H�ew���K-��1n���C]��L�p�ȶJ������^a<$uM�/࿍��6�a�m�g���(���MX�\&c���zqR����̤Q�G��&]�������ӽَ��_��:d;�)�t��+Ѣy��v?��w�� ���,wAN#g�,0O[����J���݋�-^
&��Ih�e��ڵ��L��n7@׺�a.g,�
���Y�J�Z٧�F�|w� 8�UD�ث] ]�<Dȋ�,��N�Jrd
��*��H�<ȾF�D:�Kj.��a�vqw�o�23�1�
�B��ڄ�l�����%7�%��g��0��W�A���k�G��0��o�&����8�1���l�#1�hd������U�GXb�i���
Y
"|~q�,v����A�"6A��QI��1�d���a�8+Y](�Y*�_hӀ|�kn���ЌhN^�ٲH$��A�Q5��b�R�Xg�hܿ	̄gBx����7��h�[��&��� ����4{~-�(lj���ϱ��6�Ȥ�Uh���N����.<��K���i����$A��Ɇ�2�Y��0j|N�BxeC�R�X[,�vM�
��h`�o�:t���C���u��5�����N�w�&�r6W%tߘ��5�~5��K%������r�K��8|���`|�f�bN��k��o�DȊ{7&-��1��[���ȟ���9���<�e��.hv�6��`�OY�Ŕ��1�t�^! �4����&�I��X<-1�ܩo��@e���X��+�.�ދa����*j;Y��T��:���t�jR�;>z �o�e�����.é}j��k��'�2>��`�cq�6άWgJ��V�����FP�8�)��pD��f$���G�e(*���Rf�?����l¼8�nnoH.�դ�.چ&̪9�ZS��.�x����b�;�K��HN��I"=���o���=�J�kϬ�jIW9��z�G(�7�z
(N�j5�z1OV|���X+i��1N�C���嚭�ŕRxn��%��T���$u8����O��jށ��Hb�����Q\D��.o�Q��LA],��v�n��q���*��3� ygf���+{�5�7�0����Z��􊡿�y!�|��(��*���.}N�>c�0_���T�s%���	)���֪8�X��,�%Ŷ��(+Z��%^�t�N&/��`k�X�(y(�$���>�m�XǗgP����<9w��/�f� �X�գ��W�ߤ�nn�3�M9���w��l�u� I�n��a���;M���X�|��a��{��揵TV��a!YX�%u�ʞ^1�k�S��4���^a�f������>�;�&2~�5��X�>�#y+�Y8�����1f ����S��B+{o��$�! ]��ϗ��j�\� hi��$��J[��IaU��s��9�$�Q��:#�tP[Q��鐇)�ݛ��~g��G����y�F/�����7��_��
���ނJ��gᘥ"B���e}�F+TQ�&4�Y����ut��)U��"Pb!Y��";��B�at��͵�H�GA����=~G�4=��5⇡��qk�t�+@��g��9ZAa=�	�)�n��6,1�Og��Q�t�&!�	�3֐1��(���_-�>��w�6��3�H�P7��o%�X<����.H#�	"��d}@f��^ SkM~J c���G��Sb�1z�f7F���1�ru��HA���^�Ck��3�
D�&nW�qٝ_�	w9���x�����q���`�d7)R��O\���*�R���nGb�69����AYc2C�In-gH9��꼵�q$S��K�B��b�-�@A<*�XZ�P�v�1t��@-fg���&�ɏ9�O�2XJ%���(��L^������v4��T;	~���Ns�g��^�:���3� +2��ݱK�?s,��.�/�Z��t�l}3�U~��4 �Fơv����(z�R�O|PUžr���A����.�h��j	KQ�o>0+)�����a�gV��S��u�a��Z3<���w�D  �%f��Bjq�x[��T�EXj͟Ֆ��s�!�.wV�0��C_�?l���R���LFS��/����X.XV�T���3����>�;3�G���A[��<���P~�D	B��=AXd��b�ϓko4 �~bwMbd��hS �r�qc�u@3�q�z�l+�����ZR��;�_���I'В�*�t�@@W���@������ E�ٱ/�P�"�Ğ�rx��o�.�iχ������z+
F�ɜ�պwƓ���|]�>��0u(q/��nWa%���,{9S��i�kɟ1y�t����z/��V�	5�$����7�a��1/�df;A���i��B�4܋��j�����$�;�[�ֶ��L�(+[��)�G	�!g�\+O��GV5�����%{�|������$x�4�XF�|��Z����@�ϑj�(3y�T�� N�Hz��Z�EW|6էo�]�z����q�F8U�HG�#b����O���10�����J��aV©�����-�µӲv�c��%��di{x����Y6�ɗ��.JL~��i3�	��`��_�y8[�а��A7&����1j�pX�8_�|j�|��h)���w@�ʔ'�O��Jc�A��~�+�\�p��ϵ�f�,GϬQ�o'� ���%�J4�d�������TiNu��2@�^���L)L'�'<�7*���Li.C���J���"�8���%��G��i`��z�e��$)��f^L�)�f˃9�A\G�񂚹����Y���^��r�ڂ��S{
�AF�(?�#=�{��[���H.��C/��_�`w�.�z䡾m�#�vc�t� �=������)�:�[����mHs&/v/��<ԲPɪ>�ߠ~��wZ3��FErAe��z8˚Er%߾���� ��PiBIX���t��/h#:qFi�p�w�9I�W�q�;,�t�Ì��>��FG�Q���b��1����A�6��U�d��5�M��d� g���;`PŒ!�g��~�?.�L�켭+�4[ Fj�|�[��&�
�QqM�M0���fgF�XJ���:�9�W��n�pkw
�Ʋ-�4
Ł��UŪ��j�T~X�R}ʾ6KX��Y�z�\K����TN����5s�ǳ�f���_WE�g2��u��
g����5�o�,E|���jl��+����H�kF�@���u��oGȼ!2i.��M��qI&���a� Y^W�k��_�g��� �D�!��6�GDI4��F���X�$��bg������L���N<�O�<�Ç�sH	z��7�`'�����42ǔ��qDsW����)I],��1�T���7� ��>y�z�T��a��A����PI�3BB=�1�� 3���c�1m�sQ3e����^w�hT	4���5(b6â��?kȈ�n�ڈ�̩?�d��#@��
4k��ɯY�?nK��9a��&q�}��n��	u��=�|�	x�:+�L}M~k��}�f�J��y�٤��:���@�R`+��O!#}��l��{?R��m�%[�V�g`�jl���hH�5lk�w}��jRQ���}�eAQC�h��a:Ӂ��i������E��O�֟�y��`M�q�ܾ�/��"2���������"qQv��ʴ�Fe�$�Lf�8���a��ZU�:Mx��>p���PZ������Uj�3�?@p��מ�6�����^z�Z�ĸ)f����89>t'�����'8S�d��P;	�Y�ͣ�� ]�=�<[�R@�՚�P�M��q%e�2�:�v�BN\} µU�q�2���`��Nře^;B�f�^���s&
U������b�-����܄ɯk$�R+��6qɶ=?Ԥ��q�DB�,Fd}^�k}o�)�ZB�_�B�`,<2ľ�9��	�=�>���,�33Qt � ���L��/g��#���V��N�f^�G	��w�kV_%:��S�:˅��bu=7�)n�[���ANJS�?�:q������\��ٌ���5c��h���.XnŰ�~�a�{ɘUe/J��# ��|W&�L�	8ϧ��d��C��q�6F���]!rY��<���O�l���ٳ���+ZǀD�O]�9���?��'������ 0����<0V/�'�0}�����������`�����|a)��o�h�'Dfn=UɋU�v�;О��)�/>7�c
�`�$q���[߉�����C�����T�F͌��,ZF��(RV��'[9��/:+d-��m-�w��W ؒ>�#PtK�^�|̈�c���b�*y�������]�����eNr��/���Kg-G���3�]M!�WR�k��5���^�!FD��M�yu���-�O���W�@U +<��q�̸���7d���9-OX"�+��,�������=$�/f���m��{��jJ�iU?,綟�d���~~�Y���3��R���AL.u�d.͠a��Ȅ�+�k���N�ѤV�(�D ә ��]f�;�j��^�{vݻ�fz_�0�T����%,<U�`���1���g���������a�v;6�rl�.}v�����m�JU��^�©�D�t�]W�H���%�3��AE��h%Ӕi�f�GR�e��Ч@��͠��W��"y�!R@�;HX��s�O�&�B����'^��@��`�^>�vL�C�*oa�_��]���5:��4�F��b�^�[�����;��D#R։�F����_�N_wp��~����b��{^�ѸH�G�{p^�=�]�<�A���\��6�W�±DQ�2�Ų6�*���e]Gl#w�K��X���T�/��G=پx���lA��Qɢ��C|݁�c���U��B��|	c�����_����Ch�s���J�fn�F�i.Hs H�6o�g|P%��:����o�:�B�#wO�ڬ�R�TF�G;�(����MfQb��
���Q��e!��I��s�k�B�d���^ ��E�ۗ��3�3��L�L�*��q}�1��ڢಌ�(:��*��VҹHl.�J{a��łP|�Ֆ(�t\ZH���A���}�קL���Y���3
��P{~'���'�N�;�_7$C�Y��ǉӰ��鲜��~����L�c�YP����{��$L����>`���+��h�¸�U���P��o'[��1��;t�0��d�,��ܯ�6��ZE�|����9s��ߘ!U���,E�(��흠G��2�\o@�^�Cڻ:���V���冘Kwa���9c�B�SK�_ࠞ��%ؓw���ͭ��l߿ �@u���m��8!NȢvv_\!�k�݋K����7hԧc��P�����^�����UƱ�/bo��Z������^����55�ݬ�p�G5TÁw������˭M�0��*Z ��>���{�=��p���)6�V汁M,�_>��S�JD�:�
����/�B��+�P{=3I�"����cJ׫��ⴜ�"��]A�V{�Q�l:A�T�u�L����~��-q��ñē����"SJ�*F�Qyd���V�)�4,��8�v���Y$��M!z�U��=�:��r51Y!�+FX��A]6��#���c`5S+}�g�Tq����Ff�h>L9�=4^Ԉ�ҏ`��p~;!�2��IT2�'��h���Ŕ� �����7�Zuc�9�����7��s���x�e�g��A��9�\�J��r��h�C&Y�,܊�!E)��si�ڥ�u�G�M*wn��5}����T����h�(]U|i���h��Mڢu��为��8m2r>���2�=�ԩ��P��E��T�Q����̐�qZ´�:~O�ύ����]�=M�D�#o�M@��D��PyN���:��I��]P�<ڳ2���M�L����BF#;��>0(�q��}�Z*�[Y�Y�}��<:8E͏����ݹ|�R!�S��ʢͺn��R����t�\)X���ZB[[*o��$��sO�ڀ�9�$��ak�)�`��r!���l~�e���l�m��Lτh�O΃��5��e�ב�+���_��A���n����A�XTa�@���m*�ɶ5�z���G��_�	��*�(���5|[�ġ�g�^xK5�%����R	>�x�F~��pq�J�������<��
y�� ����h+M���r6��ϪK�,d���O���W�����T =	�_�,ss7�5(��E��)b��hK���(]�B=G��\��@KwJ
۹��H�Wxq�)���'���̜��Xp���CU�6��Dt��Xe1�f"Ѩ��;��Sd����˱��-M ��5!��}Ql�_��=��P! �.��]ٵq��o��?���ϲ�zŹ���질�>��~�=����P��t2 ��-F�u���"Wa��nvSJ/���A��UV�SD�}Hl~��� ��11$͜��n7x��!�W`L#���=���)�T�=S���!����$�3B�H�^�2=���{ 8)�m.�s�3_��	E[�KLXs�dtE��@�0`�{��E�$��#}��m�E�#�6m������u~��-6^}/����M�{�C��Q�����3�T��rpP)EB�u�t'�IC�� �Y����@r��A���]� �*.AYW<��KW�j�s]��Z4�|'y�F�oc��3�h9? ��~/J!,�%+\�B]sO�ml3��q�L��_̨y�Tu�Wi`�������E�j�#W{d�f �����bʮ)ѩx[玐^��8/�� ]pg{�e��2�
W�XC��>* ��j����lR�ڐCC-4���,�%�pz�g�;�,���~���˪�8/f�����},Dk��,�2�ˋU�Q�W���!�e���?8��Nw�P�/>X� ���*�Crg�J<_T���r�Z���f�����BG`4\����q�1��?�.����t�������&hG���;�U����Q����xcU0���K�$9��������P��|Z�c*�!��<�����b.�ݴ��2�j�Ի��������(�h{��׷�!�<��7c�.�$)n�/L�-��V;�*�/��[�5��``Yk�L|��fΔ�ȅBC�1s���} T{-K��VX�>�F����H`[qC鏉}S�J����y�J��"i�@�?-1O/�$�,:�̯�J�Y��O͘�/f�2P�5A���#�[ܑ���|J��>��a���m.!�Q�h�>�lc8`h���!l}(�t��!N��A�C�&�=/F���?��!����¼c�HB���]�i?a�%����5��5+|�uMӓ/�ְ��dO�	�G��Yz�L�|E�p֌7�u������)2b�@�'J�g�'�Q��]92��Gm�
�Li�ۋ��"�&��F�l"�[3���!��	)�N�$�ot�U^�Ҟ��I�@U�[�؈cs`��S}�#�ve�KK�q��Ϣ�_�����҅��Eb�{�g�m3f�$C1�<���yh�
*ݮ�<Dd`#�Q�������+f�M,RLiSr��*턾�T�6�P-?�<���e�[�����y�c��p6�=m>�_�ؔ"kgZ���j��τ��zs�Z\�v���;�Q�4.�īGE*-\(%��}��Jgh�|g<�;����8��8%�GbS$s��A��SZ(h����0��p�&=R�2�J�:��uF:�����A^�3���Ϊ��)�4&�d6�7���V҃Ɣ���}%��5�g����j�~�p�����z�O���v����a�Qtڍڃ�F�t�9]���eGƷa�­pu�	�l�^�L��!�~`�/�������紴��+��+������!m{�8��Ϭ�r���xW��[������B+5���h���x��d4�$���gt7�5H'��䟶�tW��CR�S.7t�@����ZE�Ƽ�|%�E�%SEa���|�(�%R�,~-�VA����c�p0#O�Hvl\.�	0(��8��G@i�Ŋpâ���X�Xs��YL��>.��xe�x��"�[�ꣁ���U�/8$��n (b�Ȁ��Czy�K4nE#�9G���!?�0x���(o�o̍d3��aa���>}>��h�����2��I������
(�a���z\8�~�6�J�e.Y�}C��+��;�f�M4���9��6��\f�O���WM}S�u�����
��J�r��x
w�=_F���5PzX�h]��cn�A�n/�,� ��,VF[UxWハC5&	1�jT��H�rlO�P��.����|-���q��La����H6߰� C�?�o�pg3bf1�c��<�~�8k���mbUI���u���p�!�~�o�d��-S��8ط�8-�G��$Xl�;b��v�P�ի�1 �w	�{��f�/���}�5i�:��]���+L{�I�g!m0Qř��Y�"�K�2��aB��3pW����V� �Gӄ"�,�r�6v_mi��?�L�X�Au�_\���O���r�@����EO��Y�ؚJ����;H!����v�v��|9���E+ՙu�����X]��6�7�j�^��'n�P(�8����N>��L9��1�O	�W�t�0�	��,/� ����Ёw����k�}��\\*C���*��!����$�o��~X%��}28�w����Jv�62(�m�:�#{r�A;�:쫻#�V��"����	���<�hY;i6�$1x�gǣ���'Ҭ���3I¹R��i�y�6�j�T��-pW�Ab_��hu�筍`o�ʜ�X�A+���#i�2��ǯ=~���k۷fH6��mfL_F���ef;�3]ܖ
���&i��	|ܡ/�
/��)~V�4oz�]�#���~�H�GkW��l����"�]�Tk���ATf���?r�e! �����M���:S�CM���88���,���s𒂽���i�Jb�љ��o����X�V#lf��N$o�c�܊�օ��zp��L��F�;���tG��N�5k��A��~0�R���'l��I����6���-+��u�_ݼ�T^?S����'I�}�9���KM��a�u�������/PHzbi��v,�6
�*H!,�I���DU+1Q�Y�fZ�2�?m�Qݦ���bDGRc�n�2�8C'��U&��Kh��%�ZvNW#�v̊e)�b�l��;�\�$�W�պ���V�/���9
f+,	w"�� h��N�xt���4�ubL�N�9	��%���7��#BD#ݧRޞ�a��/���r�UQ?�{��QG: �E$� h���i�-�gYl�?�N*#p������'�>'��6�E�k6H�N5�>-4Im��ج���nY���Q��k�����vc0��k*��l��3�/U�l��Z�]�n��d��v�7���T�Ũ�n�K�T�����ٟ�C:��=)pTE��0'�������கR.�� XfS{>�4gXA+WP�5�� W����&�,�%�Ą��9��5�� n���S�C��4��x�&��m�8�+�y�C�Ly0�*'��8,t�5�(P��?>�T+�02�&b�*Kf[TF�=��-(a�s���&� ��ĐN��AAP
����ܠֵ�����(7�����$���Gv�xm0p+<�?e���$��|N���;K]S):Z�ɻٻ���f'x��ڎ!Vk�4^���yo�&�HvRJ�c#�߰6)�D4�)���i�p��'�|Z?��,u���h��]�$����"Oe��N�c`}���s��m��+"+�0�F5�0��c�
+�+���
Q����{;��A^�͂��f����"�v�ֻm��LM��k$�a�Z�=9��J�J�X���Y�;ï���3������֣�)�F��u�>�����ߑ�E���w��>73����Y+�]�D}��:���G�iy��dߦ�<A�ȻV@`�f�͠�f�3�����vq}�eCb�'���X�<?��P�❙���-B�@�+@�8s�%Ԑ�u76 ?Э�� �K�a ^��+Ñ��/5�f/���6Z7��t��kT-�ytꊹ�H�,����&V�!�z`3"!B�[�������g�5+-,V;'<�4�+��u�b�d~�(�$~�qP=��k����g��t��w�n;2i��������͖>�
e��"���#�)���B�kp��e�A牄<��1�������O���7Ř$~Sh�4�P$U��oY�<��.�&�3�C(�����Tj`���[2��%A*dIn��gЩIR��J�o����~�E��)Y�$����}�n}m�c�`�{�2��N�\��ac�#��aXH^~�B�\)����H*N�	��U۸k��?�i�x�z��(�8��������q���h���UXl3�X �-.�X�	���_�Z:u�+.W*%�]�4��z:D��D}��h�mt�'�<##��ن�9X��a<�pR���F�=N&8)�h���[F���H��(Ω>�]!Z��BQ�@7��+�X���X;�9��M���^���0�TĴ����W޳�r�D[�p R��lQ���A��L��C*
�Nz�g��(�1��H
GHO^�G1��|��ٵ@���k�y�WE}��āb�� _i<�ًW��o^u\�<){��=BM�v���-�l���B�Z�oX��zu�H~
_�ɛ��og<��)�".��s1[�ȇs��%bTK{(wf�ͮZ��i"���p: h���I�R�yކ�R��W�ۨ�Ю�c�����X��ݿ��^W崑�Bu�r�lW�k��A`:z�Z�#���l�0�.��y�Y�v���(� �Z�!���΍	��.�Ad��ҧS̩���g��ӑ�$���hu�</X{l7�R(is�+=u��k����I��`��&�\�8-��*{:/��!E�Y>6��6�Gm˂�k�}j�c`QJF���lЂ��OK0'�X�IR��a,�8I��?��K�\U�O�;�F.��X�QDTآ��7[Z���BY2Z��<�W��i�/�)r��E�B4�dt[d�򰚽�xXhpg'�=��(X���D]6����'h�k䟧;j��$Evv��C��gM!R�ClQc�����7���p���������:,��ˎ�Jp/�7Q� !�s��W�	6�:�I #��I�f�Nm�/������� �_���֖'C-�W�'Zڷ�)��T,4�6I�l�>w�]�9�a��E+C+��杗���F�MF��\"��4�FyS�ܜI��&B#%,�:�G�+E�O~����>���"�����+�n��\�X�^\�qُe[��M��I�(���c���"9ʨ�@������6��yj5)���4�������%Ds�.-�D���t�Pt���v.��:w�7�����E�&�#�	��B�G�h֣�E`[�{��D��4%���t^�	�<jN��/�jZU����.A{��\����Ն�.M�U���X�uBL)�ٛ�i��/��@V��OH@��] b܅��,M�hD0�2!vT�a�a�������E�DL�*m�{ea��K��LJ3GIjT�e7��5� /#ފH�{�;�g����8�ɤ��Zda���:sa�A�L�OP�A���`���=H�yXG��f����fxlO�N��Α`8�譍�Q9/~8�F�Y�g�r �|+k���H��Q����J8w�i���GvV0�B5�U�¸Y��KU�nA���.�"L@�r�Z��4?]44���]
;�D<A;�ŝ�g�OxO/���-˹��5�X�p��EC'�?�M ������ֽ�?�s�Ep�5�;�L��8�#����8�N��KCE����멏h0���*�-�=���L	}��3ؙ�l9�>9�,�����C�L�/^tE�.�����R�趞0UC�Ak
�?>��+���uh�W���[i֌B�䃫i\��Pe/�(�Р��OL+7����q�Y� �)�Wv(��R�|i[���UEt����;��(cK���@���i>y���S糄s�F�f�p"L?ӉQU.��Q~��	�y����� ���ةuGW�?�!��%�}|&���Y�We��0�����[H	h�b��MQ�$Cr�	�6'��jI�<#�v_���wm���(���2gd��~Ƴ�몙*\W���}�C�C���E;�#EG�ߝ����O�'J��׃n����_L�1�}N"Q��]�v"�s,�r�jm�MP��o����8N*���U\���	�JhTko���������R �Q(TD��c�:<��?�ʋ�;6`���ދ�IU)��t������f�b�17����a�[��w�:�g(Ǵc!�[�lLK1�?�x/OٺFVf�A6�(������q��d8����mJ$���d+���6v�b�F�C�M�zg=�3�8�R:ˋ5U۟�#P������Cmd l��rޯ��2�М���t/�+�s��oz޿8�r�53��+|�z����Ȇ�(ޱ�&�7n��ˆ�,C~b�{3�b�
�[b+x��ۻy�~<k�����?jLBY�r3Sw`<kG�'��Ĩ����(��5��~HzJ>\l��-kT��\17��C�����M�/��H��#�5P�sJ�����S^��
:�������>��d��Fa�f	��mcCN���,�Q���ɜ�
+�nt��E�V_�z͸� � m� #	�7S��<�� F?�{�vR
�3�",6�\�jD��y��u%�҇&]BL�%e�Y�!*n�V��:����?�<�X��i^�6�El���`T�M%�엙�Ƥ����m�o��U��¬�,/xu��"����&��ą�!P}
�����l�X���EZ�!�+���.�R�{
���e�c�(�6ÅK9,�pl�=³t��*NB*'PE�"U��'�W"�j�;�*�._$cE�݌��:y�f��5W#��i�.��M
ѱ�6��K�� gG�8Ll��C�Te�k���m�i�**��-�s�u����P���B�N��oT��s���羊;�SoD�i�[���/�Iw�: (��HT���t�"oF'����Y��\�Ecs��E��,�\�I�S���"�G�ouNs,X������ ��nΎ۞�w���n˾� �꒽kӂ��r(�:.N��6�I沣�v\@")ᚫp����`�����A�p��k6��s</E�x(�������� ��p� K܁g��o�[c��ίg�.�6Zf�<x�?�����`���^�75�{	
�=�M����O���3�!VNKM�)�ia�n�Y�+u��J���1D3��"�d�z�v�20�ڦᇯ~W��R���լ�-mH�d�7�i6h��Jx�oO)֦�Y�)�k;'#���f"���|�뽔2���r;p�_!v3)���L���t�w�I9!��xQ0爇R+��D�<���ز0��6\-c�*����K@5<�׈e����7�䠒0Gk�!#?��{R�!3b�G?6�P9=vRjkUp�\�Ea���" p�-�F� �!�.|*f��Yj�A��'N�$�>����ߙͻ,#8��h��I`d@D	X�,b����c�q��SD)j�%�;K���G�i�6�9.Ԃ!����EҭӐ'zQ p^�}=�%U΋�i��Nw���V\��?:9�a�7>���央<�]&/�Y�"�˪���M1LЁ*�Zݱ(�w|8|u�j��\W��xj�_��W!���B�d��}6�Z&tWX4������
I�3gn$�!�U�	��N� ����bz��<�Q�PQB��)�ʥQwl'n4ںTZ�<I�5+�/o����;E]�����~.�����{���~iКC�D���˾kVM/d���j��U��	?� P�u	����;�_iu��%����N �r��B���xw�@P��Ձ҃+[)D�&�B �FU!'���*�`7;�P���8�������lvi��%&�L).��T4Z��H�g�ud�:��w&���"	�0�6x�8���C��9�o9� A��G[}L�H�Z��������v�����^2?Ȫ�)#UQ�<8��ط~7�����7��G�S�n�;��A�>$��4X��ZX���0�������:����1��	�DTtR���R̀3�|E�^>P���vd�=A���Ga�����\��J̑;�l|��d��|Q���4�:�=-м����OP�|Հ�kf��˧�IgA� |�Hm@۶Im����h��Le����qҎ(;��p�q�x��[�*^m�z1�!&N��^G��c��]�K<�Ʌw�>�V�~a�;[ګG��SwNn���*�ιs�֎�X�?(4~�B�c�h�qP�� �� )6P�1�Ƽ�`�g��˥Վ2�L��a����c7��Н*�\�H���͢��^@�-�;������;>�V��
�奷�[4�"�AP��2�;)|6@t���Q$xS|1���a�2��k��� ���ت��7�O9Ɲ��9��d����������}HO[�޺#R��	D
�� 6d����|���bh�>���ռEY���U�c�%�)�	��j�����v#���_jeN���(�)'g=/0�Ҁ����`��B#�y���9NO׽��V�/L��}t8O����	WX���UzoyE�.b%�b{�����W+�ئP8�)y���%��+27�ñb������dH��hZ�D��/����o��-�d�m�g��y�fQ��h滷dѳ������]_�1����>D��]@�M�����j��X��Ϋi7W\=�0����<EͿt등��b�lE��,�c���(�.�d�=��-"���
�����u�e�N�4CX�#�bR�	(�l[��W�f�<�$��,��qA���?2x�����f:��`F[��^�����\��S�4����=l�-Rה�C�@�$�q�e �6<�>$�u̗����Cn�]��������!Ey8�%B����9�,�RZ�������-��A~H��#t�:��c�0�%�AV�)A4xR�Ԕ��kK�}��<�4a��Y(���*�R>�@l���h>�ӒY#��@�A���b�C����ç\m����;䜣����Ild�R}�B�;�'"��k.�"��I��������%+�������1�H!.���JV�9S�㘘�(e�c<�_���?�q����h��ح�tI��`o،Yx)�(ց��l�B7y�����;��}
�,g&�m�5cb��0��Zv���KW|��?^�2C~x���|b��Q�54�_�-�>H����t6V���s� �ٚ�1�w:(�3L�'5%�D�p{i�aϓ 5l��I�Iݍ�Һb�P�u��DH�:����|�~H5x�N��S��q���z��~��ڄ�g��j
uʭ`�	aF��pSJ�P��MX!�؇�^�Ua�ٳ#S��(�C�eհ� ���X-5w=Zޘ�5����������FJ|��/�7��Y��}����碦�h��A��yGw\)X�X�o�U�Y3e��C�f3D��N/����t�97�*g���0� ��j}R��Ud(T��>���E�QH�u��bȿ�"�)�uҍ�����M�"/��$P(rS����i��C���(T.�O7�t�{7�ޙ}���R��������6�e=�����Z6Sbu�k��̿nR�K���v��ŝT_R���U�P�� �g��/&D~0����g#��s���֦
�u"Mi���}�fƤ���ˡy_ۘ{8��"V09<Y~,<N:N@�KP۝[���p>��z妆-�4�m|�<�*���>����&�G��:�:�=��s���m���p0�zBGTDΔ2��O�����~e9�9�,2�� ��s�#���}~M�g���pN!�xk��mQ*��.h�-�/㎳��!"m(�����2���$��Fe�`�l��s��s�	X�J�58q-�<�	��,,���Τ��<�Z�Y���(���hj	��u�����r���0X�*��0Tj�tc�d���z�fe�z�Jj�N<����v����
���� �#��f��� �GnpM�p)O���г���:>M��4�Cm����1�..�S=����W�3ʿ���5$�_��r�"�\�!��_��[Nc) 	����rf=W��&�f�ױ�__'$�I�B�p��ӑhD�g1�z(X?���B�>�Z��Ӆb�����T(fB�iN˿�cT�fN��"]���Ӵw�n����)^�dR};�Ea�,���1��?��0^�[B�A�o���W�gȻ�Hp ѽ����A�(����� ُ2#>@!�:[�D�He�T�*X#N y,��+r's2��8sO�#	&�<z��J�OS���@8`2��P���W^   ��z��z25qC{8������}���;|��6�l��dZ)+X��YʺYi��{4�M�Kq$�0��Md��~
A:%��lד��oSF�!L^Ǳ�Ȇ|��K*�8=��wHP[+Y���U�C�:v�ک}I~#���o�>@LdR*3 x0a@(�A	�����0< '�D~�g�	��]��I��Edt�[�Z�;v�L�B�zb ��n�4�W�V��e�����9��T��ٛ�[M
��A҃����Qۡ�|�X\u���W��V.�E�/��;8G%@�i�N�pco�G��Dy q��N$
������ۘ#4?������������{�l���^c����!6tZH�8P9~p��jS�1�����k�n�ǀ�\p�$�Z�:���ׂ��aR2���a�+=�7d� 8��PD&²�ȹs�|@N��r���-����H�Y�ia�yo�<s\:c�v��L~o�Q=�x��t��c	�T�>���YU�
��#�2'&}#��D��	/���}��iN9
��@=�����B�rp�.Rqıl���-�I3�'�w/���E��}�v�|u�I��N'��nݽ1g-��.UL5�S��h����q�Y��,���v�O!Cy��{�,3rh�f �w��o���T��q�k&���Or>��("[m�ob@У����S��� ����Ot���d�k�Cww�����s���&��	AxG�(���C�9��;��"���㎢�r-����W]����������IR���/����V}��*�.=<����<��^�+���̿�ǹq�1�����J�W�˶�ۙ��-�?��Y�����}/M�)9�arwEy�����8��X>�)+�����8Q;�M����6�7��;�z��[��4Y�o�����*Y�0�����zI8 4�e���Q���	������G�} ѥ|K?�<��wHK= v�i��V$��x�!��^���>Q�PhV��?��d�E�I��*�������RP�D[�ru냯q���Q�z�8��^Cb���9C��>vc�D��U��$��q{�~f��=��ⷠ��h���L\�T����������L���֞��]q�'Z�hc�X^?� ���-Κ�k��Xs�6&�G��C��FB�/X�1煺J���!1����߯��y F�֐�X�G���\� =@v���,bZ�=�m���}�`�ncf�=�{
�yS��.i	hd�jGgV�И�%�ft�a�NU��wY������I�r���Oj$�5����E"MU�z�� p��P'v�C�y?�G�ofW�H�iՊKG�����X���\~ U��eǡ�\���Bw��p�����_av�3�^��\�Fޅ$Z�y���X�{�I ��]4������Mc�����H!%�8��_�؇��l�}@Z��v�d�p���X����$�{�AE��4�}��V��L�~�����$?|2'v�"�	m؏���:b�!��	~W�,���Z�B���[�T��Ϥ@T�a��#����D�O�7~�f��,� Y���ϋfBa(�9�p`b!�y�қ	��������O�ĝ��!ǐ���&\��S���"�뵑� 9�%��ް�Hoh�e�	��]�֗�7"��bq �P:b��bj����?�9�B�f���)*�RdB�1��!P�"��-�	��o~{��oxW)ds8���&�����1^ZH^�q�\��uS 1����#~Q�@�W�)k��&�R{��q���#]��x�<qv�6J�wE�9�\�:�?AN�Vo��	#���"�՟N=�1-ذ�_ox	�ƲQ��G����$-AN��D�L�%tj���9��u^�}oo��"uRF<o��Y���䮇�t/h�<;[/6������b\�4��+����w���p���]M��n��Sk���־�'��(�)[]���z��m]F��v� m��]Y��6�U<�/y#4�Ee�ӗ��bR�2�V՗�C�b@�u�ȯL�6<j�N--T���e<X�o)�6&k���
-�Y�@�F�_� .��ϥ7���T����}�C���]�m/5T�q ���_6���H ah�h1�� ą��~��h+�Kz�N�d�!i�L@?�9bu)�RD��=סo��qM�Ɋ�8[Bo�J!&r��WL�R���z��̰h�����|ۄ���)�e������K��BD$:���*���������6>�ڰ���vE���r�K��360�� 1+V��esl �`_,<�q2���;�x������O$�����<�$9Q� \��Fn�I�RҘt��$��҅1��r�ҏ
�s;�Ȼ����ѵ����І��90ܬZZA��V�}4��/��
���!���<�̆8y���+| FtW���f;�b�gZ�cX�w��q|�F�x�$��q^P� W�J����d4�� ���5ζ�x�1��.Z��t#E{����e�bM�v��k+���4��g�s�X�s�B�/���KJ�I��ie�/!��>cS�A��g��ZM쎭?�1���u|��]���4۝{o�J������PSRL�}���	,>	�0|��:u��C�`���y�}vG�P^�'�d��h�N�܀��Rt�h7���23S���"�"��>mn�������������Q�:�D�ԙ�/���|�	|.�ύMr��C�0{+1<.��櫺��~�� �ҪV\�P�����bT�%�F��'lu��G� ����w��h��L��Y���ζ�L�{�W����^s�����b�v߀��O}�/m�Q+o�6������|?��;��sZ�Q�T}���@�[Rp���ws��q?����ݾ�+��ȫ��?�'(�\�Y؂C��4�Q7��dFHĽ�����N1>obD+�l�v�|�!�!���	2�6����(��&xA�l�d݂r0�F4Kyb�'�Νs�����^����D=�T�Ʀi�������4���+�3�kO=8�j喕J�����������:ǘ���Ӷ����~ xvA��{�фm�H�	AX �ϓ�Z���v#��>˚������4l6(-�+���ݴ��4@)Ѩ����X'*��E���[�/���;���[,�_tD�����7Fc�,	Ʌ=/S]-�f}���?f��3n߬�o���&�q�-�[;�3;fܦ�,��:Z��{2���b���ju��a�MdB����ي���+[3i1+�&%��
ס�����Ɓ�7�P�<}i��H�e�����{�^���M�o�¦��>�gL��� ߥL�m-&� }���ޗn^�&�Rb=���Ad�_9�fզ-u�!T����r��L�L���'�0+.�*��S���5�Y�9:�\`^���5Ei<��DQe�C�J`$:D��a��Q�4$�<��'׏�`#�D]FC��Pe���Y:b��؈�Y�x��F�5��?Ǹ�1��� �ĲX2�px��3�qK�^�����.�$�3f@�f@��1��i�R}���4����0w����^��_YJ:3�N���(e~5��a\X�����]�� ��V�y�!�#��[lގk<�����BOz�eB"~N��O"*���Y����%��&�8��q���Z�(#ǈ����r��6���+{!��f�Ϡq�㸻��B�'#ڗ��v���vRI���}�������Ó5��!N�R��`����$I_����ױxu�<�) �����:xet��ٽ�X��'	�%=�C��]T���M�&œ��q��%��E���lBs
��w#%!�~�nv�H���BJS7��"����5Y��<{��AlJƸL��a��P�v�
%q�ְ������-Bfd�2����r��3�	/�Ⱦ���*�ܷ��W���>:"g���Ă���}	m�(�[e*/D���r���5Q(���n���^��I��nl�$�֐�3NO��򟿙B�QV�%fE�V4rm�����uʿ*}ٔ��W縸[�N]��H���&�|K9��F�� *�9�c (�2����fM�jD��-*:��i��t���>�k��Jk v�.¡\��1s�]l���A�zE�3�3a�<�y4���&W����� s�J����1�Y�_`n�~qD�"ݿ�#�@<�z�m��ٟ ���J;�_������=C������~ebu5x)mJsc�f���#D�"�������T� ,�r�� �7�W���c�{��؍�-���O�<�->�怋���$�����3)k%L>�_i(��"����|R��JA@ �f���7��+��Jđ;���u�_ޅ���K�w��3���ԣO��@1��ۼ�H�n*%[
����r����
�n���� �f���,V�4�l�:�o��͞r��[�IV��m�*��N^M����m�Et��Щ-wA&]���X����=DX��V(_9�<��F,{r�R[�B��$HK��Rϳ&WW+o�M�A��kP�+�-H�u�)�>@-Ӗ�Y ��xz஦�^��@/�)�qN��M;#԰J[)#^�/��F�%Y�p��Be�|<�<U��s�7���e���_L�7�Dk�s�2��<"]䝕��$��\���om�[P�"b�@��m+(fڤ^��.	�"�e�ʌ5���X*��n�5w�Д��8C^�~F�ڴ���{��%v^����/I#z)�M�t���Qa ��=���m�!�s9J��ul'ET(��L�^u# �$��^�8��Ʀ�� ���d��U�i�U��/���[}_����߼�Е���$�|Iz:S����M�
h�[���x�V�XI�G.8��X���`'WWWMY����O�I��+�&��re!A���ɜ�$KW� �m�h����Y�&@�+W<�y��J�o�T�Α�%4r���u��c��O�Fu,�_u`���*�Ā7���� yϚ��s���A�8��O��F(VlZ��f�?bb��gb+д�˫��^�S�j���6�]'�/�w^ձ�v���!��}���J+�;~	����&Q}o[ ��˵�1:ƨ�d�����iaZ}`E��v�l=!'��	N�~\0���y�I�l�� lx�u�<>���{ng?>�����ģ�K��TѠ�'�N��u�ZCF��kX�����^Gb�T�j��v)�jA�q�J��63��<<�����֠�4)�嘺�;D�+f��鋻�(��DQM�.����#؇��b�t���L�	�ۦ���q�b���������%)�#|�'����>;1���Դ�9��Թ���/����i���Hr���s�o1w��C|�pE
���#�� �w�-⬓j�^���.�ٶ a6���%�),=k�����Q¾�G�K��8��)�eZ�+�2�v�R@
�P�`�����e!7�K+�Q�F>�
 �#fhɻ/�s2��B�(B�\9�b�<����Y�mie�;5о�n�Jty4�0�G���4u��YwAGD� ܆���hu���v[�TA��6��F�Qt��t�#ߖ(^��,BP'�K�
�4��%?��I�����U�����9BU0#�p�&�)���"�{�q��N~��`�A�ȝ���ypK^&��A�*�H���F.V4�.Y�RK�Ή1�o�+6ZQΠ��m�+�cڻl�|����f;���i����Hd*C�U����ldO�
~��՘�4,%�N $:�f[��֮)On41�.u�V�P#0)#3�)tB���jq�t��I���-��<wN�0�b=Ƒv���f�Y�l���)*�(Z^���\�e⨱(h6y��Ps1���ӠF�#��̷D6����B�����=�"^����z�<�iU�S5D!��xݎR�r�WE�9�L���O�KX/��1gv��F%�y[���A֕u
��j��3x4v���a厍�0A[C�d��ړێZ���Vq��^_(&�Y��������a��ɂ�fF0�9ΐ`W` B���<��)K� ���k�C�=QO����:�</��#J�M��r�
����d�����|�!T���`l��Kg6��N����D|�Ā��K�$�;������HHz�0Z�`)t�-_ɩS6��x�}Vm�*���yݲ�aR��LL8n��g����JܛJ�X��)��d�xi�����$���)?�r:���?gu�^^��ssʚ.�~���y�h[c���!�]�X(��)�(A�3�M�w���"\���a(nx:�Jc��<²����_S'x�џ2_@�O&��S���|}�tn��1@qT�F�D�:�����xL\��ܖt(f���rldG����[L��T�IK��r��Yo��A��20q�:mӷ�O>�J<��cTK]��Mmt�)����Ku�-J�a(pץf�6���e.].�Ԍ��i��S�و���t,�X%� F��3�*�v���jd��cvP+�|�sb�ch7���J���3}GI@���ݲ>���)�O����O�t��,s��Q��K�v��./5��|��9�需���f��k 7(h#����6xw��zj���`s��K��sA}3 �C�u��N�h��&?�~� �p� ��qy�b(@�,b��'f���/Jq���*C�1s+�e9�}��ɛ\d����{}>�.$GWk�!�ٹ�i�������d0���V�N�O08��[�� �����c�Ї��Vکڤߕ�a{F��:�HԽ���3*���r��x:�����N��g���1��f��-�����6	�����-�1E�7�������K%��?�'��=����>��<IZ��ɂ��TVV�P�֡�I��z�e��L�2|��C�Z�x������,T2]	��2��x���NgVs�G��[؉y�vhsZ��6TD[5!ǿ���		��u�n*�dsw���ID�_�������:�يMYQ��P��3��mH;~�Jkt&ee{�Խ_m.�~���
��w�{��l'zm�=���v�ɪ��׷K3�-Rd��&����>�j'��Y+�g]���׮W�f��]��5��n��g��o���7�s<��h�$��}}2�/ȻU�">O}�=q�J������9��a?�r�]t<�K�-��_����y���|v�ww�e~TE�׆�&����ʓ�6��gʓ�F�`��K5Ο�Ԭ��P�]�_Wn*D���r���z�Nj|���p�-�-X
�h"g*!�n��\��O�{6Ϫ.��b	���H����M��(NY�����M��$5
�,?��,�S[XrR��l�R�u��z�)sC��lB��@nҺ�M%�ۗ�~?��l�kUys�?Ғ�(�X��d�쾼qY�B�L'�ϥ��=�����ܐ;��wS�D{���v(��{X�%�sP�=n���;G��C0K�����dK�^����K��b�ys�^7�"G�ilC��mj��0��|��v|���Zr��f�ۨ����{�����=Ej�70�,��#��EO��r���R;�D#�����ʚ��!4���6��uߣ����e�h�Ymu���h���=�g)��?�-P۽�	�9g�H�J��Ԋ���8�A��q�ʋ4*�bʻ(�\9�}k�?��j���o�imjqG��[�ǣa���X@�/���K���s D�Y�0���m�?���fl�8&�5�T��+t�<�Ȃ��'��K�'GS���q�ŷ��$�_�)�F7Ұ}���3S���`m�̚V��p��#b]���@A��z�I!*���D�TZ�\��̌��֌����'z�4�a��iS��)���E2e�2�����I�X�$/43��t�3�Z�b$�<my��?{���C��K�~R5��'t��N��(�CdV��Ȓ��;��0c�߶�������[��jd���6�������H�3����G���~���ӝ�`����>+5X��O�^�[�< {�Nk}�[T"A�%8��@ �K��ԕ�[�����x8�n�MР�D���鎒1�fnDZ�:I�t:�F..�"ԡ �|Z'S�S(��"�����5�3o)	��>����� zQd�U���`N4{�"���7���r���;�&�)�y�}�ϘfS�/z��j��6�� �8R����cM2�;Լ���W���B^�</7>�g)���r��c}ʖ�Tu$ެ�v�/sv%�h�j
������ ��q�ZPQ�϶Tb��k���5鋽�%�ʨAywq��(l��9\��Ő�H��:�J�Ppj�&��1$�I��m���/�e��+�� �Q~��Т���R��`6SV1�ßV�y'����P�`�����0��j����4��]}�/�=q1K�ԡ��{��5��3�Y�x?�F|�d���{7��|b��ʏ̹y0"�~������Y��>Z~��M���fT��hZh�'��G�� ��Ho��a U��1�+j�Ζ؛n�����ԠJ��zV�T�;y����e̸��9�2n�O����N���?���g���Sr0�Dt�H�Ƕ�#6��e���g�\g���!�w̽[� �ힱL��/[c �J�ר���5�:Ȕj7'�u������ ������Y~'���c���
j=k�ߊζ#���3*�P�;�(3���
	� Iu�iI��-,�BJ?ɹ���n���E1�"R��?����h�-D�L��w����� b�#rJ�49�4���$.�֗�+�_���.:Z?e,����,&W��-����-У��� �`���6 Q���}��B��8be��h�w��O(�(-$fHig���-5� �����������$	��VNb!]d�*������]t�qf�K����� z�T���O��y7�p��Y\`{�k}�.���Ѩ�P��x9@@BzA ��"�S����Z|�.!�0D���x��NH���}a�QG��T���Ĉ=$�B*�+���� � kt�K��Y�fn��F{,��Ō�y�'�����r����x:Қ��O����m��F�D��e�w��#r���t�N�U���^Vhϑ��������k�26uG^4SJ݀4�tB8�b��*�b�)�V���/&�F�S���ir9)aΒ�TL�1�_��5���%�a�;��EA��b.�H��4yɨ?w��p�K����)�rلXD�oL�B�$�9�m�_����g	�6����E�^�0�_��4m��='�/dK�^����d�lpʟ�$WM�棕:�(R�P˼�C]�׈��o��!��g�bCZT��]�,������.��眓+�]�?c��h*1zZ9��X���g߹}^Ch�*v���X>�<ݭj/OW7�@��K�#l�H�uґ,�4Y�d�)��-�IN���v�U�g�/r|lɄУ�KG�j���Y\�R�\z������r1O/G|�e��Va�RB0����P���Ms��4���Έ�%9`�|x���f�������dN�gCj����4�ʠ�jx�� ��p�}A�%\�~�n���^�pi͛m�=����(�
/P�F3�&)S�:���^{?��唩8[�����n>�����ɥٕ�]<��%�uc��r��0��A��y��.c�呸��
=�4���<i�f�Bf�Z ��+e2L�羘́���t�`ՖE���@�A^"�@���g?ߵ�<���`obT���uc���%�����U�#����\�Y|զ*� ���x9�}�3���铧�\��n>�3�f�3^XE������L���T��xjS��L��R%FO��j�dwT�u�F��������fX΃y��v-"�m{>��l��0q�f��@:k�O�����q:�d�Q?�Ym6ݥԚN�Y̕ϴ[�Ŀ������Jla̈́�u�u��_�rxY��=Sҹ�	�sTɥJl���&Q�����" �{��3HaBP���c����J2��8���^�5��q����>Խ|WKշ[�b���5\`�߭{�6�S���c׃��(���)%s�E�����!��;3~��+m��)(V����o{� ���)�0�(�9ۺp�hF����`��vE�s� 8mπc}Y�۟6���l��Ȃ�r��I�Io�R��Y�&3����t=#A��t�#�������4feR�aݥ�V����ϣ�]ڳܡ&6��ߖ�<x^S?i�֕�_7�@�MU�H>B����3[g	
��ci��H���X/S�)��GSP[a����M����%L��(mQ���կ�鎊�d�L��ž�Ik���A8��6�0��:d�{�"�;2�B�J�Z�-'���d�$?.��ǢEPUw��X��/^�6Z�.��U�
�S?~�}|gZ>��a�܂.Z�2��w��e�W?PM=Bb+��iԜ�#Z�_B��nI&�=XL��SL�Ŋ:B��λ���u�(��.���~Nv7H�$=�^L5���zi!�e%����{���]�k������P븀�ޞzz�9up���j���On힠w�k�`+O��4f�d�nK�_�E����)L����X�����^2�z(�b��|�٪����Z�P��Ъ��a��U��إ�ڧ�qraO�tw�Q�l���E���>�,�Sg-E����P����'~�W�?��/��d
a������r��L��M��]pa�e�����|���z;!�t�"jZ1�u�����֏��3K�k����ǵ��t7�,�wǽ=y��c
�z?tX^��`����z������aR}�L:�~�m�����Y��Ť��}��R�儖seY$�b'Q,��[� 2���g��M��W2���l�i���kpSt����z�B�a�W/2�	���a�2�u��_^|\��n`xu�mg2Z�
Bl� e~��,q�I�2������x�:�I�bâ';���i�j��J��[��l���$#���b엑�}�D=Gʢ�VJ1y��В'o��9�k�2��Y�Y�ڶ���貏�|#��Zf=�)��\�.��}��]X_
?��ݝ����`p��v��e,�Y��g�kk�9�?��8�"`�I�˂Z���㹲���m�V#-s�]� �/E���~Y���"'E�B#)�F"P�a���N�����Q���g�G�ͳ��#�r��h���ؼ�ł��ܤK������9&�z��%�[��_�O��&����y'|���E�X�&Ņ<<c��#��IG�=� ��Z/`y�i&ٞ"-J;�
�aM���'����k����?�/�����1�kk��I1��[� ��Ȁk
�ӑ�eq��2J��O'�q�s��	�Go]�f�n�����X��N���`)�0����b�!�$듨N�r���K[gK�7r%��D�T1�*o�]|�7�<:�K�STxH���J��;�M#NQȄ�v=��\]��s�h�oM�h�����p��4�7�����W��'jG�!fv�+n�yٯ}�
��*�b��Ձ�XI�����D��գh�"�^��������##�E����$���F�f�I��{e=���552�s�0fp�fZ���S�1��u3����l��m���Qc� ��y����̿P�F����lk�����&9h;[�o" �|F�m�T�I�w_���j|��Ӯʈ�}2�C���Ხī;E$���x�P��wG�]���b��ێ6`2?�$+����AJ�>��k"�Td�C�*\*��"��(������<��+��;�b�BLoߜ�"���(>�j�{`*��)R�����u�ȷ�i/�*=���Y�7û"������I��2c�Dݹ���.��*�ZfH^?��(�
���,�"_;|;�;�v�y��Q�Q��O8��pB���ͺ��!�`��竎`F��J����/��3ӿ��;ٌ��
�@I {�XŦ!�����#*�IςQk�\=�L^�Q�T���}7��
�{�)V��1K��5��pg��<�i3�HK����c}�*qZ`�H�<˅���d�>��D������a����uӎkA:}�js}��O�X�r��8�Rݵ.��sY�J���-�� Fu�_�[��
�cz}��U�)$�ʷ
48��=^sܴ�Rl&_�<c������+x�C�M9�����\(�#�ڒs+��_�2*'�������Gd�LŹS��|�x֙�i��kì�������T�!��:����<�O\d��:k�)O���]�n���ڥ��hÃ�)0�
u=�E�vt�nm�Q���1�'�q����rA�~�j�0�"U��{������?oe����f|Rq}
}:{U������ٖ1"�w6��a"��̦��B3�_�~�$�����cLu�~?}�3�1��I�l����N�Xfw�t�cd�k�oC�̈�\� ���|�o~�h��	�Xũ�mW�{؉�dI�ڽǂUl��RȧXfW�������E����S/���.��n�&�Fv�����s��;�,�),�)�$Q��Tx�.5.�ʿ�C���P=M����up��p�!�#�C 7�E�J0Qq�\��4\m��
K����Q��i>�?4��z�e,fs@Wo�&�O!j�P�x��X��
�!����]!	V��ʆb����4�d���1�^n�Bdu��?�,�F"�O�����*SX�m��I,�o��*�4Ӹ�T"��~\xJ���K�:A��q"5O�J��&�J��+{�7pEpz+���N[k�E�,bOV�Ub7y�SS7u\��V��l���z��=�D�ɋ5���x� ����t�2�W��k����UG|����u!�d`T?�)���{�B�i�uծ�R������=��2����%�k^jqAθy�ޖ��׺4�^��3?��<q^PK_�����D�9��۲~׳�B�x�M�Bp��;�{hY�����Lq80s~~=Xk�o�	�a�����^�Ԓ��l���"h�a�BGq��@����?�����z)�,��uδ�	tsZ*�_u`pӜ���L�i�qX�O�����o�oD��%���[��x�T�~��x�h8[�A�~ƹ?lR��"g*����itn��^F����8j�8���{�#��B&-��)6���?<c�� @�]er�\Ĵ�S��h�@)��o�J��zJ&�fZ*���F?��Ə��o�0��I���Z��#N#�
�U0&����/����ߪZP2Dy1��4]�iM�o�,Y�k/}7SCf\X������y.$y?v�r�:����+'p�G�D�Ή���96�r��4o���Բ�'qY].gc�JO�e��(4󐍽5e��N��E����,u���U��~�$m��%��D%�k��ؾ%�nF�0�C��х4��jx��[������vX�8K��C����ɃUr��ǲ���bue&#F�W�!$cܸ�Pʮ�e'�0�$w{��.ܒ���e��!���_�v�^� $��km��6�.�b�A!�Fɑ�>x�`3q�q�e���vJ��֎6�ۙ<�����E��7�����%�$c�*yr�29�M+�5��6�҇Z�h}(�Y'7�"B�{�v��e�O��I�6O���-��ҡ�+���5�:E�L�����=c��V��0��Z�|ؒ����2X�ϟQ�,��>6#��	���m�^]��Ŧ�[��s�ǳ�,�ku�5���3�=Q�iĘ��CR�~j���֘��w;���&������9��?>l�!���kH�:�.�T,�Z�͑^ݔ���Kjyԥv�z�~[����쌡Q����s����S��K#2J�����ޑ'&����F�6'�g�L��_�(m��H���e�g=�C=;H�/q�l0+_�{�<��`IjK��U-?��:,#681�̴����rS9^��I�='��!�A���f=N1�_�t@ B�@?�߭*K"g�3~�#~xћ�\rd!�v4=4����C��-�#JZ ?W!Vx�+�5�1t�nw�8ţ[y���<5q��/���"TR��oKUH���t��	M��0Gk&��<`iF����{q��������;�����CIY�4��=(>�:S~(P4c�#@8݋��{���Z`�J������g���s0`X2s�T75C�P ��+�c��%(��8����?[��ܐ��]�Y�7X��ã;I*vfe�
[x0H٩��S�=M���-��B���Zp�K���f7�B	���>U_6�+�+^�� ,��ŕ%�m��D���{ު��,`�5��Ƙ�6�/���*�I�B�O��^���.��@��憩�s��Wu�H�vg;��_s��B��T��7X�/�[��M`��?�<�����U���S���&��t$�F��雞��K2;I�|�*ՒktL���N�I �۞/(�!x���bEk�XG����� ��������!Ӷ�|ؔ�<�~���VCO:A�5j�_��ڡ7 �u�dP�1����k<Vro!^푖���`����ç
�W�Ǣ�X��:�*>���2�F��?:�����@�5���G�Z�'g�ƘKs�哲3=���k-�IiARz���!t>����/~�>_�\�^)�6v��0�R��2�l�1O}ث���8�_9I��,�]���'_̭ {�pY��|��Z����� o�P#̈��W�T�.א<���Ξ��8�l�c5(n��#��|]���T>�!�;��7��x��������o	p�@IV�e�P��k.�/@�=T�C¸�C1WEٽ�5�rZI�~�@,��c��uvTt$��`�~
��L����d�] �G���	iy�F)�O�xT�%_l����~��'��1BͻY�j�^�9M��e�J�r���D?��"�&KXl�=��@<�{J9���z/�$X��?ub�ƻ=Q�䴒$�����4�[{�� M D�h�U�M�'�bӊ��A�So ����u���Ð@l�V���&-��(?aF-�~�&�|6���g�M�ۂ�f�L��H=��he�g>rUcq�qϖ�X����7̸�;�/;Oew
�Ģ-�^N��'Qi��%��{���L��BFZ�k�T��#�TN��A-��V�@�+����PR�E��X(��ٿ��$;l6�2�����'$��K�me���ğ���`�YYU��&6�3�ស�@P`�,Ƶ6� &����[��p/�/��V? �B�IgD{6>PZ�k���lb���c�-֜�(�^HR5�3��Z��Q�ٛ��e�"�A��OC�0,8[��9G�58Дht����mNj��D���v4����)�!�䆈���ѣ�#F9u]��V����"{�h�ʃ/_G7g`в`Ei���U_`_|��l�6�M��Y���<��+U߸4�j��x�=�Gr{b�:UG>��E��Lx�QN���ƥ:� A�����D&JS� FZ�=��-ᭋ�:P%��d�-�r�ɉ9�u^�t�q�!�0�
k ��3S$��)/�P��	�	�B��:�%S�G�1���O��V������[W(S�ʓ���M"��qǈ"r�Qe���A�1F��|�kQs�Ƣ`D�� �3z^�뢆�|�o�?��ԟh�K3Ǽ~��)�d$;�L�v���ݛ�PʛJ"��±��ϐu���Vץ�W"�B81���[!�+/�3T,Aؒ�wU�b4�=l��F�޷s��Dq��hV��V�ُ2'��3-�Jf~OA�u ��S���%�>`���z�\�R@��=����?n����o���h2t�t��66�}���yR%�].ؓ�sPP�w�L�B���yEBvU ;n�WyV��Т�u����F�:��%~Df7Rw�Ic���Q�@j���egV�|�������읩�pٵV����~��bUɶm.���S�}�{�}bM���c���/a��Z�1�LquD2�4�M�e'��Ku^�ߖ�i�'�)���<��k�ṛ��X?ʟ&]���"� ��e{�Q�w��ɼ-�m�⸡UV����`N̰vz�&ee������j�԰��u{�?˅���LKw�YK�����c�{(�D����0(@dNO���ɓ�L-3��6P�c�Q��C$��J�Ee�b��ѥ`���fp��_�2��I�_�­�FCE8��V�i� ��qY�C{�%aW��.�AZ.~{jWP�9�ϙ�`~z]�b�����X�Q��i#=~>1�15;��JrCR��[�M��(��̒�;��ٺT��{���ӂ~)5�Nކ� ��E< `�I�*�H���ۨ6�o��B83�yN��p�3�i5�����=�!<?���(Q����a؞OP>E	B"��6Ԇ:a�H訾��1����ܫ�mV�Xp��El67dXD����i��(�L���̲6�Λ�	�1����Ar8�(����]�� ����(.?�� �.2E�9�U�9o;�N�Ç���0)7(�.���� �	�]!��j��dh2#N������s���}3��8�Hħ ����l���sK���}�D-#J�f���P����u�rH���"�(J��k���fFD�77��F��_k^���t�����K�.h�p�6N�� -�dp��RZ�r��L_��S%�<�&Yͬ��e�r�}���A#��d�̛����������X�����Y�Ɛs�ٹ���z+�� ��M�6C��td$85([�v:Z�R�����O^�@�q���{�- ���쁋@/@>_��#�x'q���ү��6�&�9��f�6�s�5����Z�
%�&�qo�C�;Xf.�!�m��,5�6,���)U����<e�xt�Q��\�]Y�{Z�J���դ��r �]�6E�M��:�
A{7�.(�7'f+��	E;ں{G��߷&5�A6�9!]���d��l}	��f�>^�{l�D4�y�"w���vZխh�צ���{�#�eD=�3��Yڟ8�(O�3�nWs������b�sІ�4���)���ʚS�w�\�ҏ��=�+�����h�WUN�1�-~��I��n�Z�j�>��0+,$ �4��ޓ��>��������l՗v�j�4R���g�0PqƼ�?���:����2��w�P`.���Ԋg1��I�/��c}`,<4Z�_5OV���+�dj='ϵ�-�����IoX)=*��`E` �6ƀ�V���f�Ƴm9**Y��Ҋ��a�U42�d2/�jΎ�0	��>T�Cd��,�..L�0�mbn�}3�%�i��?O���L5Oh��`�(@�\�dWZw�P�a!�`@�A�p����o��_���<��-�����@�:а2�о<X#�-�G�����m�N����3ǉ��X{����O��K�W��>A'��oT�Ct���[�E���,dk?!.��4�O{���U��G2���`Ө�m���2y�J��u=Á��o��=n�v�.����_q3�7��/O]�2��(����u*=[FD����6�h��(�>�7yAz��X��A��YW�"�sOYQ4�)1ԑ���.$B�ɠS.��i���&9����x�MAo�:�9wUe����ML��x�K�]�q��[?�4\�X������گ`_�ƾ�F<��q,�q V��X�ȅ�a�#>��]ۇoJW@0ZA1���g�����~�r[t��)�����]�s-����N�xF�Ț�{>�ü�Xhm�.y�'��N&~�)���F�eK�<R�&�~�OT,ZGS����2�X�~A���6�� �$Y $��wi�Z	B�/���u��,C.�{���� 0�̍M��#�]����s���Jn�x�4����F���d=���y#�����i.����^x tv�;6�z�^
f� /��u�����=��@ǻ�XÐ�ygH�Rur�����a�myu���u�~�rBzvg���1��P,NB�~�b�N2���v/�Q1SZ�$�D�֬���z�U�ݨ�����ei��>.�X��p���x�������Sb�d���$M�6������:+E_v���<�M� +��穞p�1����'��ݷ��weB���UcM���@;T�Wd<��>z�{�G�G#��4�H�@ �O�v�A�@B��%�i���,��E@����Ľ��S�c��IU�_��ѱ��v=�Y\����/�'�0s 5 �����:�WSI9�BRZ�Jf*2G�PA��yh���mR�����=�5>V�յ��Amd���H���!�N��k:Pյ���j�-�f�J��B�g?s�|��	��Ҍ���d�F�;<ל��v2���9��-�%��P��<
�o��Pf~�\`~Ch�b*%���\k4�bG?$���ѥ�_�
�~_��.<M�;��)�ԋ�ľ���cxҋ$���!ldj��6a�"��y�C-�U�3��_�=�K�(;?�?�IKuaq��x��A�H�6�'�֬�*�ƴ��ɚ�}j"%��L����dq�e�X�M��u?3�}v:�ozMu��w�"J�=<�؆��t���p�P�S}[�m���S�ޮd ̑56��c;����ވ�G�=ѳ�p�+V�sp�6�O�ځ�5^��:��
$2��ŰnxF[Y�(d0�Ξ���b�n����'0o�~��ɵ�Y���)��,�h�7,��	��^� �tK���wΥ���>D���U�H�5=>$_/DH*�ĳ�\M�&M�*�#�:�J`\ 9��ɥ�,������0�[�M,7��tRE2��U�4�ٜ7&����ƲSR�7Q�xZ��'��n��P�߈lB�犄��f�ؕ��S~�.5<zᷦ�y�fv$K8(�������f)و��r����8}�'ׯM���%��3��	��0~���ٺ�'S'�H�H:��S�{����F�ҭ��K~V3^�19��$ތ������h;�yg��# �]��8yK'W�~z�ŗR�v��>�n��|�j�읻u_$��E�u�G�ш�;�N-
�[�DV���S�S՗�]�%{p�[�t#駔�k���>�����{-���?�V甥�S\����6��-��.�E?����lWxDkf��C���K,wSik"�>�`�z��l��RAV��;0
�^-��A�+Ԩ�߭�o��wUc���ʳ2�YD�������w�'��&�c�V�^��j�1�dl��uc�Z2��+��T
(����x��:�4S�lQ�yVPװ���)(qoG� k,�Ņ�D!���=�[U>�B���8`����x�%_�ܼ�!m������r?r;�9�*�(C����rB]?� v�B�Ѹ�"�5��0y�xF�N"��p�,#�`Y�w�܅"�Ǥ���Fx�-x��
(`c�Os4�dE���dP�RK"&v�6S�R��@����F��	P�8풊;�F�����߻]s�T��`ޜSHS�x�J����a�E����T��~��Fq���aK
��=#:n���r땞_��M/r-S)��+�����{I����f��L�gbi}eߜ8�Dq� �{/��t��'얦0�i���$Fђ�@���z�O&x�)�kj|=�ú�։�y��wA&���#��9��(� �����I��W){H;�4��%�۞}[a6���,��E�Š���7�浔TЧNώ׉+6��k>�2��?e��	�a����ڒ���˷3{��Y�K�����Բ݉�N(m����S�K&���=�>F���mN����mS+]����O�O%Ώ���9��U�(�A���,ƞ�{�lYe������c���BPᏧ���9��C��6���\����VXh'<�	/Xi�e�Ea 	�/��фX��3���s��u=��i���J�K9�[��S�,����4	ٷj�nIeh����8m�`L����)�s���H�Z��@�1�Q�ʷ��d~�w��!x �ы�V��Ô��5ʻ��J�:,��V����Q�A��y�О��%;�8�e[o���ͬ���E�c�����f�P�#���s�y��kr�����׆�n�9O�M*?mΥ��F6���*�0��E1��x���	�m�N���Y6yj��Vlq��@����xr&u���0J��=���听�*".���)���,z	�~�'\�b9"_Wq�͈�s����G�l����T%')�s�>��mx�;���O���^��h�0�	�7��J#M��P�a�� +��;�t+Ye��]�gz�����,)��PY����-��7����5=xOާ�s��	6��.8����?��m���e�7i�p#Ǌ^(�2����s�T��|y��t�Q��`����t�����T��/{��w��1�6����4����K*kS�"�.Ca"2����?ܤ��(�.DEX��c?�L�G�x���Jo�0�k����1���,k�f�2F��D�y'}��!�_��m8�r�����8��w��l8.Wlm�e��-̆ �8��ٚ�MТ��B��e�c$?�7d�S��CN�۵�
�c��C�Nc����h1�O���F���(Q�>�Ī��f� ��Q� �pŢo8gu��c��$��dl	�����g��o��MV�.��lku�&�9+?H�; a���#a�L�r��`L��4F�̃G\�{Q�z��Y�n�
�+��u�e��_'��ȓ���v+��G�h ��9D:1�/̢�C�h��'Ŀ/���\o;E6ųMM91r.��_줄����rْHᅹ3����֪�����xK�km���#`E�t��*o1
GX>���&���!��E7љ ��p�]w����C|���f�#lI�	I0ȷ����x'�aڻ?���Y@�[��g�f��x}� �:�5g��2�\�y�߇��YJ�������o�d(������k^ ?vГ���+8p���S&*�aR#�L�H����>w��afI΍[�<�M	�ƙF��s��(�T��0ٖ:�#���$ֽ�EP�Am�C����޼��l�S�I�_�\�?ZڃQQ���,��Z�'n?�[�In2�@�³��A�N��}�Nd���s#�b�fٛB����7��+x������2>�	9�����	��`�)pv�05r/�Ϳ#[M���{c�0�G��q���R1�B�p�W����\�T�k�#���8<�.��,��R��F7)�h��dH�d]3yW5�Z���PӐ$��O�¯}k2��TK9SP�9�w�r[^�uR���O�"��HW�Co�?��L[V�"qꂼ��zǞ����3p��x�#��fF��%����P���3	�$xVI$(# ��)���h=%�R�Ҝ�?����v�Nw?���3.QNw��"m�}�n�����{�<.� ���'l��V���
VΒ�ͭZV?d��o�m � �g��\�b������q��>nOzPU�k;���˲�7�
D4���)\��vp,��T���?�,ڔ%�t%���ek���$�.�P��|�~L��?pj�CC���cMZO��Wn8v������Čγ��ѐ�͂0�Y���YЏ��
�����#�t�lC�{���ܪ�NNz�!��/�Z:�>���x�EA���K��J͊Z�*<ɗ�=zd*2��`�G�DVJm���W������h#B�E惕�|j���6�9깩���sT�}}�h���՘�}sQ*U^����Q�@/f}�R�	��WX�WLb~��ݓU ��*�U�Q]�A�3z�m�t����������y ��E�H���Q��@�Ϫ�w�1��J���!_48B[���g���ݒ��
<�y_�iL�אY��Ԇ2��_����X�CqT�� D�[-9�(��O�f�ȳ΋|U�RLj�kL_��+7O73o���di�LU�8v��DئT^b�O" �b|)'C5mf��,l\��w�"@y+�j
� � ���ĺ%Zag��Bo�BC��K������Ơ�b������W��5F�pC+�D%�`�q�~�o\��h|�� M���2ݲ�D�x�� 0�y	��R	����\�݆��{*Pww��������!�!3�wS�y��J1�2�7�	��Mb�E8�"Ǫ�4!E�"`+�F;��ćb�x�� ����A*�<�W��{@	�+p� �'��� �%�eAߐ�>r��ѳQ�~O��`�l6��1� <)�[��;.�B0Wv��?r���D [GB��NL����޲<Y�'���n�ܓ~:�ȼϚ��<��H�w�/J$�oM���A��T|�prD>nƿ���ay�Qim�{�'M#]=aF�t�7jk(�ףZ��@{���B?j�
�ۺ�e���i�wq��x�\k?����<���
@��)��6^��^`�zc>$�0uN�̨�J#��љ��`���b�`V�)��F��g*Y���8��CaVo| ÊL�[c�87��ff�J��������+��Ld#hl�m�[Zfu"+�-ɴ�s����<�d�GN��v-'9n�*�ÛE���[�x�<7�l -'������Q�v�"-�:W&���pW�e��)6��?�K�䥔��X�np!�Ї
��ڭ]u���I�!-�C�ˤ9�"�z�cV ���fúǫ�32�ŉ���\�:C$z��YLŰk�.0l����L�뼝Dv����P�OU�E��je���/��γ�X����pKޭ��,���S���xZ$��0.G�=���i�0�	&��W���s�a�S�)��y"M�L~Ĝ%�D��6�́	{��ٲ�p^����-�_7O��݄E,׈uu�n(�k���>;{��H�UN�G^�[M�WsY9����%c$S��{j-tP
+F���*V�L?Å�.�N���Vr�vz)x>Ěi�V��&�>W@��9K���w��E.�Q2΁�S��p}��V05�V�2��a�d��v�?��Q��R�0PZB�#ʉ_  <�x@��,�FNb�o�����p�n����K�Tq?���i�q�fPʓST)��Z�k����yml�J&�����b�x%q��*���lgFd��)�z���ޤ��G�_�@��Y��I;�ŝ9u��3+�B@�ݡ�O��lzJCt7N0��,�g*R=� JE��no�!�gTm�(����A��]k��l�Z#�ԥB���C���>�
��O>L����<�Y+:�o�`9/&�K,C)��-���l�R��;7-�.^c&��|��iC��z5�(5A���~�H���N�m�S�$vIP����5k4no���W�ic��h�32�o�hK�ԝ%��xG�p�"u��p?+w����'�ͻ�ˑ��''!�c���ޭ)����Nԅ"�Sd�#�#">>c�t�kͼ��GI�T�7!7��Żo�/5;�^(K2[#�e)Р�ܰ�ǩ�>�x��=�9��%U�K�� )��Y�~R��"洨Y�\#��c���Z-H*�c:_$������o쩪�S$�IK)+�����NP�>���< ���.9��{�W�T�S�fVGSB��[g�Cn��Ɔ�x�,=Op������`H�O�{&+/*�8n���/�;�^��r���m�U>JI�;-����v��F���(q��D�;}6.��:�v;�5�����k�8�_(���|)(Co�Rkn�m��|I��M(�u龥���[��7#:�IE)Ϸ����3����H�D�y0D�f���Q!�T M澢��X��&�r����ڝ�c�t���eD�3e�H��o� 濩�C61�d�`%��,X@vL���1c�k|��t���Uy�B\sRhk���Z��SRF���>�jhi��)��$Vqֈ�� h:�NK�����r�c�At�=�����X�j�b�z�=�CXܵ��P�;`�����9q-���-�5�R3�/�HGdU�:������%K}#Ņ�i9��U绷+þ��S7������Y�2Z���v6v]����I��� <^�b9��RQ��Ӳ�>��Q�E�P �y����_K�t���FЯ�Qwq��4����ʝ��R��._D�s����I�p���VI�ԁX��ICW`ms��x� �:q@�}���Y����m���I�/.~)&��$�n���r&�_:"�HF�U�*m0)S�d*��պԂ�r��Iu���"��,��du�S� ��/�L�-)_w�J�ďR�a�"`7��Ǥ��;�nB�si�X!�?$�|v?�R<\�%7�a�J������g��qݑ�2B.E����K�0����X��j��ŹӬJ�Rc�g�S����.�d��J�� ���Y]^O���c���"oYn���7���1�P�i���T,)皼�v��ta��P�w1�Tߚ�C$��x`=SV��z��	3b�۳���Baaȋ����&�i�z�;����� � !Y+�L�Q�+��ik:�f�pAj���P	���A�KĪ�lB����i�oI#��������k����Էs?�L�r��j�s3�����r�9j�I�L8�+��>_�-�O4_�����r��C����ޯ��(���
����.�yTre>*-VW c�%�	��$$e/��MLx��T������+ku�3w�Gc%_�0HII��W���%D߂�X
����@z�6#�Ʉ[�`o�qO����f_�#�bMVu��	��Gú����P�����T�C�n��.I�7�b������מl�\�kVwK�^�}�:1V�UJ;
�"z0R���#�x�8� c:_Œ�����KƊIK����'sl���|v�y�ۍ�"���۵�y<��M����,/?*{L�K����{���3�Ȟ�^}˼Y9��Oh����t�O?T#k*�3���C\x�L�Jw�.�w�	6[���V�Z��.{!� ֊�3��R=���0YQé�&���Js�J�#��+M��"aa ��a�V"W��K�	�K�5z��V�ͭ�im�m��Q��8\J�IWO�yZ�=C��CS�k���l{}���-ޝ]N-A��1�]�s��o�A>-I�$�U�ӭ{w �]��˂̵��� h����t��ҧ Δzh�������Hp�K6/|,|`��t�T�����y�hU��� b̔�p��z��j�y%>����l���\�Ñ^�*�&��6z����Mp���_�	Yě$�=���#>�}4���]j�-"��+�0���:����`pw?|�o�>!V�N�q��Eto�R�aA��#7ؿ6��W��'"8j�~C����ε�����p�g󇛚�۶>�3(�)�LC4���b|�I�����5��,���
t��į� ��������@>)AY�o;��`��k�0��b��y#��@�"<�4�U:ƓR,�/�9�T�����s���B�X<͈��X�� {:r���i�Z�⹑����)F�I�r�M����2��]�>өwTf�'`�ej��N��7t�,���Jk�ZM�"�X�@��W������,7\A0�v_iu �}���ޫ���[9>��Ey�!D��\�B�����ܕL�Ό��&�uG�'k��'#�pʴ��+��d
!��X��J�A6�*Ny�vNi����α+߇�������pi�Vl!*�B���x�����Rj�rg����Qx�/�;�8p�p{o=ſ#Á$�Yr��g�ɚv���l6pW�){�>V<Q0(@���"+�B+�À�8*�R��e�&�hm�a ��yZC?��ƃ�-�g�}S{����	�LZ�8po< uzWr�/֗n&~ѷ���
D�+��
�JfOd���V�RĘH� s#����_�	7�#'��w��V<��	�!Ku$���&�Q�2|-�C�.)@���JP�h96(x15����i�����\�����?԰^�x�O�'�*l�@߆��-7�tTu@�W��݃�6y���
��/u��Ј۱c��\οi@�l[��C� ~
3��Vg�y��9c&���3G(�_��jdx�ш��Ac��ϥ����-�ɦK��G��R;��v�k9�e��fW�UPA��K����K��?�q��� ��SCB�ƕ����F�D�\�M`U�K�>D_���G�?�����]5]�&�A@���tc�����-~OAރ�_�o	�U+�k�%�T���T9dF)�ߡ�%,�֏���H�O���|��N�'�d���ח�i�E�bY)��5��!��[�l썒�?��?D�������
�¨�Le��h��>ca��'�[�=YxQ�����>Qte{�q�d�o�*1�_�i*4���+��G%���Tׅ�&��+.4^��
_*�?o��@�1��5hhX��"ڀ�qE��E���*�T�TVn�qĊ��'�9�>�BX�`�Պ�~&D��nB TZj��)є���<X@tol�n��S�C	�r���l���֭�$�mYt���2Z���~����r��޳�Z��>�˻ߤ�Kzߛ�,~�;�Û�	^�p�8���$�O�P�3��Ǔ�V�.��5���@a�����͗�0�a<�E%]ʠ(?%|3;����`ҟ�x���G��
�C���=fH����g�^��&7(��2�b��^�VRLK_e2y��a���W����u�{��x��M�Ci� ��W��@J�ݿ�n�y�=�/9#69Nj#O��ac p�_�8G�V:��c<��>�p���m�*���O5t�VYrn���5`�W��
�_��5��>�;�?���CF��]
�D���v�$M��]k{X��E�V�2,+ꮟ�F���95��M�Y��E�K ��P�xeZ�����]�_�f�A��/�m�/A����L��iJ>�a-�z�7& t�3�I�v*��zy�tZ���g�
����&"t�D��>o���x�?�ƗS�8�2'l���
 �a�nE˰7�W󲠉L���!O1�����s/���N�o�d�L�	��H�x4!Y�y�C��&��%*s�}��!Ճ"{q}���إB�;�7'̀0DzQ�Qm�J����4���:��P�)Dr��0�MQ��$S켉�]��	�6�����nsC���ô�/� 7�`7�J;J��[e����FNԒ��/�&�c�1b�?;���⸍p����+PP�-�΃U{�ѵ=����r�9��Pn�h�}{��:�ܚ�$�6�{�$�g0J��Y V ����	^_9R�a��{9P�W��O9CP��)�W���������}�_��b�����:j��T�/� )���O��ˀ����ۿ��KJ���>gB� c�	fd��'���!�o��ښ��yBj"��XK�H��y�%ř�T~����կ��4���������$�=z0��4���_ņ��y~U�����`���7 fJ��YJ�`�`R��@Q�t��#-����{;���f��nM�u�G�S�=Kg��������Q����gzA�Oi��uU���r,�m������7S�$3,�	��V�v�vs�=��ߵ,�+�����d����f
m���?)��T�A�|�zCL�GG��r�{L��i&?�?�N��(]T�2Ϙ�vϭp`�!4V�� ��V��A��2X<��h���E��h9���0��Cy�z8\ x^q�T�n���Ҳ}a.�w�vC|0{Jw�Z�~O��Usa"��K�8�**�p���E�vK��I����S��~o3i΁=��m2����Ny�c�VP�+l�����G�c�sΒ�C
Da�̍��@�/��6���q;��p���%&�ˋ��X��Jo��'
�'�+-�Vs[����Ժҍ*2�-��S<G�rj��|�D��2  ���V��#��2%R�n�w���0�eƻ�a#�Z�����!��1-�n��{�_]G�j{g�1���RKe��F���$�ȺȷJ��(���f���twN"R�KϘ�VQ=�񚜮`Y�DK�4�/�({ (��R�w�V�;B%�>���Ѯ�r~!,"�}�>r�\�ѓ��.	���q��a�H�V��<���HYCn31 5	�/�5��V*��� �G>{�� �"ہ]+��W �_�j�Ū����5��b@��5��K�?@�@��:/�u�(. (i�`��KK-D��3h\Q\�+����!�.G*;6prQ��z����,��*��)  N�V��xonzI��,LsU��R��
�OO<{�6VgwO!^
.Q���P�\_+���8��Ś�V�H������:=wç��y���sl�����ԑ#	���Ex��7W�P��[Oj��cj�*�*�GB\�u[�*�~5,�K���y`�0;�J��l�q�'�(�"���Q����
)��<L�z����fys+�L��7�I��.��EG��� �ZK�4��������\N-j��:V�?M�r 5m�sՅ�>?�����dw��w�J��Y\�r��)�&�Jzrf���	O U����ʾJ��o4�w�S��i�3 l�� �x�[F.�0�O!��vi�Tո֌�`�C��� ���3���7xh��z��)���Ufm��u�ڵm-� [8���K� t?���u��	T�)K���fv{�:�C�<D�ֿ�UH)�T�p,JN*�=┏0`��:f���k�h '<~M�V�����fn��7Fh��2��f�D�^��=���4>>EPe�C���8�B��W�{�R����W ~�(����R��5M���K�C����q�ޯ�m[�u��W&�����"�B��fw��[2d_�:LG�� "�S)�̷Eں�dY7"e�r�E�ŲTh,jsk�����
Į%���+n���k%gY0�)�7�C� �!��7R堵�����Mz�;@�i2+�d>���`�B�o�ߡ���a���_ZR��J%V��m{��--�7��Akb��8�+�c�f�On=� �`.�D�$B��R�0�!�2�n�9B��)[�LxBÃ��Z.Lfֽ�-@m�� �7>��g�{���k�-��y9+�[%��p7&��`�8<�o��=�}>F������?]��l�O����k:c���5��c��b�;�L���@�~�I=� �:�=��9!�҇�b�����p�@6+��i͸�~�	�T�a8�����,�犇D\���r�߻��A���E+������T�N7�Y���|�CƢ2�kĝ�����d׼� C����w�Ƥ�F$���1�e��_�"a����|��� ـ; �6����wP�Z&�:c��\�n��ΰ�:c�dk�Z��1M�A�V+����(0�oLW�~��L��}��������|���`߈���nY��;�h�eb-�r[����,���8���w4�?�S܇tr��\�R���v,����}�T*0�v"cp�: b�Ӿ����ܟx���Q�!���;&��Ƹ�̝��:��ğ^~�G��sS����rzK�WUZ��Ͷ���X�o��V-[�n�#	!��pE�I	b�[}f2�4��?��iӒ�U�����̚�s�\��A� �$�J�(������h���SU���߻�@۪�cy���k�h���{+���HS�1���*�7��"9��>��؊alx������A���6����4.&�R��5����x��0�����jh��`�7��A����~�Xoa+u��u9݇��QL��%��I�8p
��jI�Y�	��0��YH
��7��|.�QXQ2[-��,P5"N�'k��~R��Y�~��E���|�v��C��B�bJY���dd0���l��GG��	�r
���v,� ��O��m�*�v����YvN9�z묵�!W܅����������ې��M$7>��s�|�D]���w*h�4�QW�����uz�f0����9&2�#�N�27���j� ��a!V�7�~S�D������޽�ʓ��2��;O��|{�x��x�d�wr�qe�����ݿ��pdX�Kޢ��}X�ڪW�b'�T9=��^h٠��f�g�&�tcZ���L~�T7���9�9�B�~��.�� V�7��p�ӛ����®���k��e3m�\a=֗���N�J�����у�sREt}���Vw��k��3rn�]����v��=�aW��'�.Wh�L�f�Lܮ�D����8�y����t��� d�����1��L���rGLP����.��B�����ԱH� ����\s���cq%�N�i��|I|�ʐ"#wV#�����*�d�Q�Hvm�@����a޲�*����G����w����l����{5�V�?�^�M�L9����Q˰&�x�\���/k'���{��<?Ci\Y��9�i$���ݑ��!Gjq�I'R��7��*g�*��mĢ(�{ǔ�+Z��Q�ǒ�O����:%9.�رͺ0�S_qnqv����ѵ��T��pT+ң���(���)�X����^�Ԭvȃ	p!��T���Sc���Tlч0>
H���d����1�F�ٱt{��Al,bPe�����3�A��A��� {��s������]�܊[_��ڛ������Uؙ>hJen,Bf��"ax�ҍ��-�J�d+� �i���"�!µXm6�����(�o��_쪗��� {ؑ���n��]�9�R�C��92N��� ��myd��(���`���o�Ŝ��oG_4O(�B<�L�A��!�4�Y�J�/C���@�r70K9�ZI���{��m���c$��S�S3���nsZ��r3鼳��WXz�
�o�V�J��*���.<ǎڵOlN[v���e�8H�X���<�Dg����2�u���:3 	��zh�+���v;���D�9H"���e��4`R@�`�����	<�0�ފ�]i�B����\X��yj��9wjdƴ<�Б��/r�ʄx�1R�k���لR(����_�ZČE����a��X�,�ji|-��!�>#C�9e��S���|�
ӥ_O ��n�;ɶڌAv.�填�ʱ73@�C��˸1ђ�'�1LR:Ӎ���UCU�0���Fc�L)>�Ʀ��0�/sh0�$�r�S½
	b�6������t�O��8��"�����8��.�[eu�� �+��7�fK�i���Ζ�C����j�����/�k��1��myc�Z����*�:�o���cFZ�ns!N�fU�����֗���G��F��%hX#T�c��ǌ���\Ǚ�Au���#�������Ԣ�t��q�-8&��ۥ�'rQ�0&;��P���~v�$kċ�	�c�����=��E������(�QɽyTr�����|�;�<$1�T#�a�]���W�ͺ��]TU���=ݕT8f� R��J��1.q�h�%*9����\o��p���#��E��0l�ܖv�����.Y<N�e"�D�a�WE�Fp]) �ᚫ�����V��A�L^��H|x�9��J�*���7?��[�67��Z�bL�k=�E�4	-�W�؄�z�BV�?w�rE���5m��C��2�?���F�RAX��m]WAp6��R�ذ�c.=�����P�k}ޣ�e�};�ә���q:�!kqpR;�!ʯ��K�c@(8.24�;��_����v�<������N���'���~�/��m\JF>��#�5ǋWt��	��Q��L�Cjo	�'!W������``�mԉ�����͈'!}*D<a�}�����������7|��&MS}4h�*��o�/��mP��{/CX�[��PZ�����cR�
�C��s��+��׆����������E��(��h䧜UZ0d���3/��p|�X 6��Ye}p�c�����~�L�M�Od�ud�q��S5�[e�e�e =�� ��T���Ó�X]��d^�)o�y��W+k��[� ��HPD�ы���z��,?�V~�L<˷c�F۱-��af�Hm[o���=E�5��{PI؁X*Z���v���o��ƅ9��cj�˩�މh'�v�\< �^Y���l���l��8.�)�g���=�������NKD��YJ(o%>+^
�/GI��N�����x����ז=�K*�w����֣�������c��Aϱ�r0<q^�T����t� C�F%�AJ�Z>�]���t�A@�~I`�m�g�xt^;n� ��� a��o�t���T�Y�N{����BFX��HR^��\�߳l���p���� I�}�?3Ȇ3X?� r`(K�xz�6h7��l�$U:�
E ׬4�RcЍl�65Q���� c�V�x�]#�%В�/�TaΙC�n����vPص���ס%͔�J4F����K�2��/��,�@a0��xsmׄ*m�7K`�hH�&izV��/�2�7�P���h��3Zb/ 7��]I�;��[bB`mYu�YHi��Ͱ�j� Ԭ Y��UTd�y��<l��*sm%a��6q�ƱȮ빗��vfZ�ŧ;林��}�͏7D��`�?;Q��ǻ���R�ѣ����h��vۻ ���+C��Ы�A�[݅����N�������n�.���AOF��Q�yҶ.��>{�}8�l����Pv�Iu���A���(yu�ZE�'��b2�� ���' zU
�u|����#C>�,��1�X����6s��6c$G�Y�� ��d!�k�}������}|���q�
�/�=V������<�Մ�u��!�:"l2���
l�-���v�fҧ�ŧ���/�p:!��0%A���z$�RO,���������AL��46��Z;���QD��vXYόv�����&���`��~�e�!�N5=cS���㺻��]r�~E3ߐm"�(+��Y^�{%�����L	� h�+���$�Y�C������A;[���.rѭ�p��
}=1�g�	�WFT������2�3ST��T_�,�nO��{�������t��'�w�^�P�ec{�ֹ;�8�AU�
a�G6[��"5��u�4�:�|��Z]FH$�H�7�U�v�M�6O����;��U2���9�.�栉��jR������eUUd�|�u���:�;�*�-����]�98�ɕW���ql2�	��-]1/�XLJq��EGs��.����1��B�8�T[j8vb���9��U�)c�ؓ������f�y*��쁦G+�tjF�b�+N�fsB±v`��(v�p����)��^.w���]Q_��p!Ќ䑨�4Ш��1������,&`�ǒ�Zy��$��k�q�ִ3N�?�lHC��{
��:�qѦ���/�4�k(YW���Ѩ�����",`�Q`�}��;Åe�%�N�Kb��4,]-���~;��A�HK��r��&��0�������H�4�Ad�Hä}���$��`]7դ��^��a��G)�cO�:$�Jl�!�P0��rT}��vޡ���NH�T�	Ba�RXwZ#Y�S��:%Ԝ�a%Z"��7�Q�J�۽�Me�O�-;I�0:��q�Nw�S3��~ڜm�砌��"��@d��_���yM'���Bc=7iűC�M����jͷ���\&Ѷ�T�ް��_F��R�Ex]9�S���=�Ap���+�%?��ߜ(�e���6�I`p��G i���:�7X�g>��q����F)⣈�#����|��4�,�>M݃���#4i�ܸՀ�p���=)V�z-/��K��AN�W���"G׎�������6���g�:�NK��@J���n�������]�"��|��� c�U��}Rh�8Fx]~��Q�D�|<-x��?g����Ψi�{"l���z ���kG�y,rFߴ��5��3�����ǜA Z�d+X�N�TNA~&џ�>�/�{B�1�:���E�w`�N���-jPT�Qɵ/񒷰�+��4z��n��pX�[���N���NP@c0X\���<s<����0W^����N�.�\���S�~?|��g�F�Q˒��[��&�?�7�(�q�$� ��#$���O�4@�eCM���9���lQ�/�N,]�>|�=u\�����a��D}��J4ڄo����߃['w������p�i�T��݅O��dL@��?�)e�Nu.��؄�IR���CG{
�+-�����`��JZ���j���� �"\�]�&/���n'��`��q�:�t�Opy�ۮh56_������؊�ڵA͹ro����k����� ;�٠ú��0{��!B�d!a��ws궚�fA�����3a�)N -FP�	)ϩWg�Q*E��*ypF*+w�ys>��Zw<[f�s�|���6'�<����,0SB�R!+
@�����h��u���fG��M*/ #7l�uU+��$`�#/}��U���Dѿ>%'�o�++�=+�ml���+D�=ηC�֫���lO>��4{��}�4w�\�:�LܾP���+y	W�p!� ���=��z� ��#"�n������p��������G��e���>U��(�Tt�dn��D~Q�BȆ?�)����LF�*Yf�͚-X�Mp=ǖ�Y��Ȱ�Ѽ��H(��Xz�:x��;�<�n�+�����Jd���@��щd6w= �62�}�{����2!����D8?R�8��V�'��������T�5go�bPc/�sHJh��}�w�>�3���F��|����9`L����/�}?f�f����{����
��ز� ��4���eS�$���|e�X�D�lJɉ�	�u����]��W������K�$~7g?�9�Ř�3��C�� �q|�@"ߟAĐπk�iU�KAx 呿���P&^�������t:Y�)}�F�:��^k~Hr%z�����wy:�b$T�ܶ���p l�ǭ3���ةN���1"�p��gJ�%<���aw������O�:����.а���%�X��C+ޠ�蜇m��h��w�y���O�GK�u�t Ч�g�-<��oEu�M�΢�ڊz%uci�J+�����<J�Ik��7�ƚ#�K�����@R����3ޖ�C�Kq����Yn͹����?�Za#y�1���S���N1{{�S��A�o�8^Ǎ��D�ҝ��cL����L�9Lgx$CE��(�Y�*�����o�S��m���*~�ʥ��k!����H@"s����x�aHA���%�3�lX3T- Ys�m��mc8;�\Ⱦ�ʱC�����!-�$��4��6)қ�T�	�6��e�?O�?d6��O@��^adɁQU]�,1�MH�R����#�T��^�x�4Ir8�J��-@�S��f��CR�΀iDaz��Kg�p��������ȎC����/�����mV�k`T4��"�"�����[��I��e7�ü)�)���}c;L �BI��ܔ��5�v>}W@���V^m��X)	������u�Dw�͠��p�����՛��#�e,���EI�J�i���YaVhߖ�~�ǃ	��?0���	k��r��Z�}ᛨnC�Cl���n�`��kc*K��i��.	�1ֲ���D�1���:BaSw����Ruî�v�������B\�b�Y�����Pu�L4�a9Oz�h{�/Pg^�|
rO�L�����2E��(^�8"��(�M��;�U�3�hL�V����A�2S����y��g��/�<'`s��^]s�_Zt�AU�*� ���K�	g�+l1�C�5����
J\�|4�8 3�MFig�
���Jq�C���hs���QH{6�cO��u]&� @P������?�V�G�����/
>bGX,r�C�Aʽ�X|�,"�qw��*AS�_9�����|	J��׊����v�'խ�c�|zx#b�=e���ؽ?L�-`��&Z�2��"�L�G�w���� 7�`j��*� kڧn<����K��Y:���u��,xޖ�^kU{ S*�/�$:���*�֐S����y�izy�D3�X���	Ix�A������͞c���Nt3�E�"s��$l7�j�_�ˑ��8l���1u���6���GM=��L�:�F��y#ϙ��;����&+�Ñ�#��:Ned<$��?�ٗ��zu�&bZ�;K�a�n��������b�}%�u�i��eSxA��[Ck���&��bOv����6�����:������b����t�		Z���O�SwU+-��glíd>S�
��]���}Ԡ�T��`�wN�"���rN�"���I8k�a�/��q�y�(�DC���o9��{M��2�\h<�-���Θ��ښ�lxl� �[ȗg7�:Y$�r@��SD-�D��|��@CzX��"�!��Ա�[k����iM�oEȒ��ߗ�96��6���,��|'����VV��;ÌTk�	M��J|���\��R������0��m�-�@��j(�u�>�J�eʵ&��9�&l;ط���2\,��s�R�Î=5��(?���85��{"A}��-�$VZUP�카P8�V%�G�ti�#�ؑ�a���w�J��m��X^in԰��m�eU�v�:{aOlE�&{�*3��l3V˶?��J����C���0�(=啌X��^q�����# �I���j�0a�50{b.��B�\A}�1B`��U�j=���Eo䆒����\�7�?R9*�;�!#v+�P,��}� K�>9�Ì�6rʨ�����m��4u�~�|�_W�����p:큱�4�_��>��z��\���dW��~ bK���_*�Ʒ��q���G�2�x
��f�`�aU9;eV��-c��i,�@���NEZ�8>�:K�"�i\���Rhm�c	^���{"�U�Y�.��M�V���Bd��$��������R_c,�-L$����*�_ z��3�I�K�9�Ac�b��j��+n�U�۪���-��\ ^|�d)�,"'l����$u:�"�0�7x�Ԓ"�`ړY�ݶ���.}�<'I��]�3|Vj؝�e~������ѽV��Pi�)��X�a���7^�`��S�5x�)s�1�t��U�5����_��a��ue�H�.;k8#�X/޽�_;!�/U'ťl�p������N����{����T����\�� !��a�H�����{�k8��yΊZm��VW�v�a�l���&{i�K�ŁJ�%m?C���^��;�[5���׬.��!�ss�Lt\�[Z�@=�8�%a�G�~O����/��V��ٓ�Q�l��Mn'�;td|��If܎�*��	��*=� ��
��l�v:�v��i�S5��TF�y�p�F�1�v����wW�Pn�������.Gru��>++��B�9���0�y��GU����&���xg*5<�;6i�7��[3���`���$����4�VsO>�B����B�"ɼa+�r��O��c/ u�M(�2���Wmº��ץ�mN�?\!�O�Xx�S�շe*h޹��N��C5�C-�WZ����K�t�����½c��{tsV8�����p��������/�%VK��Ek�u(L�0�4Gvɘ�2�C�$V9ч����k>8n�規�T�1(Ğ�z�������Ii�P?�X3���~K��G��F��cjeO;��ԑ�p	V��u�)1�* [@�ӝTl@��萭b������:��ټmI�;���M�I��E�Ou��]��}���5	�}
�U��;��6�l$�MN��_�$e��}e!3�܆��VMƥg!S�v��=ɷ�2u{����f�������I����q���i}I-��������p�gf�ť"����8�����vfid����_�����C+�uK�@����!] ��&�J.�u�"n+`:��Cщӏ_Ӏ������_����ܷs��J/YlE�V�-0O����V[i�zy.c���l�*�!aK���H§��m0o��Xb���̄&P�뇆�:G)�࢏''�d�_�cX)��tQPI
{� ����i>��;J�L8甀a{F�������X<��L�9Û�ť�ѷn�dB)��-G�hx���)9�n�g� ������؉$�����t�es���[Qm�r��!|5:Xp^"$!���P���_���U��U�j��N����f���?<�|�6��)Ű���<�l4�_\�j�O!!�KT����.��d�x�g�Aq��y��`ޚ������v";��Ҏ�x�Y����H��ލׯ�~e7��n5�t����� �}��/�ci�,7��x-:VB'�����6K�KM��[�[���pp�c�ڇx�t	o���>�X&�z}�<�)9���?w�P���f��Ll}J7`l`��GY�J�wc�)�